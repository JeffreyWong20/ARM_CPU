
module main (
	clk,
	v$INPUT_183_out0,
	v$SHIFTNUMBER_186_out0);
input clk;
input  [21:0] v$INPUT_183_out0;
output  [4:0] v$SHIFTNUMBER_186_out0;
reg  [20:0] v$REG1_103_out0 = 21'h0;
reg  [21:0] v$REG2_315_out0 = 22'h0;
wire  [10:0] v$_64_out0;
wire  [11:0] v$_329_out0;
wire  [12:0] v$INPUT_190_out0;
wire  [12:0] v$NOTUSE1_102_out0;
wire  [12:0] v$OUTPUTSHIFT_320_out0;
wire  [12:0] v$OUTPUT_117_out0;
wire  [12:0] v$_152_out0;
wire  [12:0] v$_157_out1;
wire  [12:0] v$_47_out0;
wire  [1:0] v$_0_out0;
wire  [1:0] v$_109_out0;
wire  [1:0] v$_1_out0;
wire  [1:0] v$_22_out0;
wire  [1:0] v$_23_out0;
wire  [1:0] v$_296_out0;
wire  [1:0] v$_297_out0;
wire  [1:0] v$_30_out0;
wire  [1:0] v$_319_out0;
wire  [1:0] v$_31_out0;
wire  [1:0] v$_71_out0;
wire  [20:0] v$OUTPUT_316_out0;
wire  [20:0] v$_127_out0;
wire  [20:0] v$_51_out0;
wire  [2:0] v$_196_out0;
wire  [2:0] v$_82_out0;
wire  [2:0] v$_83_out0;
wire  [3:0] v$C10_125_out0;
wire  [3:0] v$C11_208_out0;
wire  [3:0] v$C12_146_out0;
wire  [3:0] v$C13_90_out0;
wire  [3:0] v$C14_168_out0;
wire  [3:0] v$C1_145_out0;
wire  [3:0] v$C2_283_out0;
wire  [3:0] v$C3_328_out0;
wire  [3:0] v$C4_68_out0;
wire  [3:0] v$C5_284_out0;
wire  [3:0] v$C6_298_out0;
wire  [3:0] v$C7_123_out0;
wire  [3:0] v$C8_161_out0;
wire  [3:0] v$C9_171_out0;
wire  [3:0] v$MUX10_45_out0;
wire  [3:0] v$MUX11_122_out0;
wire  [3:0] v$MUX12_251_out0;
wire  [3:0] v$MUX13_57_out0;
wire  [3:0] v$MUX1_179_out0;
wire  [3:0] v$MUX2_69_out0;
wire  [3:0] v$MUX3_184_out0;
wire  [3:0] v$MUX4_50_out0;
wire  [3:0] v$MUX5_110_out0;
wire  [3:0] v$MUX6_194_out0;
wire  [3:0] v$MUX7_38_out0;
wire  [3:0] v$MUX8_150_out0;
wire  [3:0] v$MUX9_222_out0;
wire  [3:0] v$NOTUSE_159_out0;
wire  [3:0] v$SHIFTNUMBER_20_out0;
wire  [3:0] v$_195_out0;
wire  [3:0] v$_234_out0;
wire  [3:0] v$_237_out0;
wire  [3:0] v$_238_out0;
wire  [3:0] v$_65_out0;
wire  [3:0] v$_66_out0;
wire  [4:0] v$C10_239_out0;
wire  [4:0] v$C11_263_out0;
wire  [4:0] v$C12_92_out0;
wire  [4:0] v$C13_326_out0;
wire  [4:0] v$C14_43_out0;
wire  [4:0] v$C15_135_out0;
wire  [4:0] v$C16_27_out0;
wire  [4:0] v$C17_75_out0;
wire  [4:0] v$C18_250_out0;
wire  [4:0] v$C19_330_out0;
wire  [4:0] v$C1_276_out0;
wire  [4:0] v$C20_95_out0;
wire  [4:0] v$C21_324_out0;
wire  [4:0] v$C22_25_out0;
wire  [4:0] v$C28_67_out0;
wire  [4:0] v$C30_274_out0;
wire  [4:0] v$C31_229_out0;
wire  [4:0] v$C3_93_out0;
wire  [4:0] v$C4_203_out0;
wire  [4:0] v$C6_4_out0;
wire  [4:0] v$C8_189_out0;
wire  [4:0] v$MUX11_314_out0;
wire  [4:0] v$MUX12_304_out0;
wire  [4:0] v$MUX13_113_out0;
wire  [4:0] v$MUX14_198_out0;
wire  [4:0] v$MUX15_96_out0;
wire  [4:0] v$MUX16_264_out0;
wire  [4:0] v$MUX17_209_out0;
wire  [4:0] v$MUX18_332_out0;
wire  [4:0] v$MUX19_137_out0;
wire  [4:0] v$MUX1_33_out0;
wire  [4:0] v$MUX20_268_out0;
wire  [4:0] v$MUX21_256_out0;
wire  [4:0] v$MUX22_333_out0;
wire  [4:0] v$MUX25_322_out0;
wire  [4:0] v$MUX28_53_out0;
wire  [4:0] v$MUX2_327_out0;
wire  [4:0] v$MUX31_104_out0;
wire  [4:0] v$MUX4_331_out0;
wire  [4:0] v$MUX6_204_out0;
wire  [4:0] v$MUX7_48_out0;
wire  [4:0] v$MUX8_265_out0;
wire  [4:0] v$_235_out0;
wire  [4:0] v$_236_out0;
wire  [4:0] v$_281_out0;
wire  [4:0] v$_282_out0;
wire  [5:0] v$_86_out0;
wire  [5:0] v$_87_out0;
wire  [6:0] v$_10_out0;
wire  [6:0] v$_9_out0;
wire  [7:0] v$INPUT_191_out0;
wire  [7:0] v$NOTUSE2_241_out0;
wire  [7:0] v$OUTPUTSHIFT_321_out0;
wire  [7:0] v$OUTPUT_118_out0;
wire  [7:0] v$_149_out0;
wire  [7:0] v$_153_out0;
wire  [7:0] v$_157_out0;
wire  [7:0] v$_210_out0;
wire  [7:0] v$_211_out0;
wire  [8:0] v$_6_out0;
wire  [9:0] v$_89_out0;
wire v$0_108_out0;
wire v$0_277_out0;
wire v$0_278_out0;
wire v$10_114_out0;
wire v$10_39_out0;
wire v$11_275_out0;
wire v$11_313_out0;
wire v$12_188_out0;
wire v$12_325_out0;
wire v$13_80_out0;
wire v$14_136_out0;
wire v$15_16_out0;
wire v$16_116_out0;
wire v$17_24_out0;
wire v$18_8_out0;
wire v$19_34_out0;
wire v$1_121_out0;
wire v$1_219_out0;
wire v$1_220_out0;
wire v$20_244_out0;
wire v$2_177_out0;
wire v$2_178_out0;
wire v$2_97_out0;
wire v$3_291_out0;
wire v$3_292_out0;
wire v$3_62_out0;
wire v$4_5_out0;
wire v$4_84_out0;
wire v$4_85_out0;
wire v$5_270_out0;
wire v$5_271_out0;
wire v$5_49_out0;
wire v$6_227_out0;
wire v$6_228_out0;
wire v$6_44_out0;
wire v$7_308_out0;
wire v$7_309_out0;
wire v$7_70_out0;
wire v$8_126_out0;
wire v$8_185_out0;
wire v$9_160_out0;
wire v$9_176_out0;
wire v$G17_72_out0;
wire v$G18_130_out0;
wire v$G19_52_out0;
wire v$G20_19_out0;
wire v$G21_115_out0;
wire v$G22_207_out0;
wire v$G23_100_out0;
wire v$G24_164_out0;
wire v$G26_54_out0;
wire v$G39_91_out0;
wire v$G40_142_out0;
wire v$G41_98_out0;
wire v$G41_99_out0;
wire v$G42_165_out0;
wire v$G43_155_out0;
wire v$G43_156_out0;
wire v$G44_200_out0;
wire v$G44_201_out0;
wire v$G45_169_out0;
wire v$G45_170_out0;
wire v$G46_41_out0;
wire v$G46_42_out0;
wire v$G47_279_out0;
wire v$G47_280_out0;
wire v$G48_166_out0;
wire v$G48_167_out0;
wire v$G49_216_out0;
wire v$G49_217_out0;
wire v$G50_13_out0;
wire v$G50_14_out0;
wire v$G51_232_out0;
wire v$G51_233_out0;
wire v$G52_17_out0;
wire v$G52_18_out0;
wire v$G53_143_out0;
wire v$G53_144_out0;
wire v$G54_128_out0;
wire v$G54_129_out0;
wire v$G55_213_out0;
wire v$G55_214_out0;
wire v$G56_174_out0;
wire v$G56_175_out0;
wire v$G57_301_out0;
wire v$G57_302_out0;
wire v$G58_287_out0;
wire v$G58_288_out0;
wire v$G60_334_out0;
wire v$G60_335_out0;
wire v$G61_257_out0;
wire v$G61_258_out0;
wire v$G62_305_out0;
wire v$G62_306_out0;
wire v$G63_55_out0;
wire v$G63_56_out0;
wire v$G64_162_out0;
wire v$G64_163_out0;
wire v$G65_7_out0;
wire v$G66_40_out0;
wire v$G6_212_out0;
wire v$MSB_303_out0;
wire v$SEL10_215_out0;
wire v$SEL11_158_out0;
wire v$SEL12_249_out0;
wire v$SEL12_81_out0;
wire v$SEL13_223_out0;
wire v$SEL13_224_out0;
wire v$SEL13_252_out0;
wire v$SEL14_77_out0;
wire v$SEL14_78_out0;
wire v$SEL15_28_out0;
wire v$SEL15_29_out0;
wire v$SEL15_307_out0;
wire v$SEL16_266_out0;
wire v$SEL16_267_out0;
wire v$SEL16_79_out0;
wire v$SEL17_259_out0;
wire v$SEL17_260_out0;
wire v$SEL18_221_out0;
wire v$SEL18_2_out0;
wire v$SEL18_3_out0;
wire v$SEL19_202_out0;
wire v$SEL1_151_out0;
wire v$SEL1_294_out0;
wire v$SEL20_140_out0;
wire v$SEL20_141_out0;
wire v$SEL21_133_out0;
wire v$SEL21_134_out0;
wire v$SEL22_88_out0;
wire v$SEL24_299_out0;
wire v$SEL25_269_out0;
wire v$SEL26_197_out0;
wire v$SEL2_154_out0;
wire v$SEL3_295_out0;
wire v$SEL4_317_out0;
wire v$SEL5_124_out0;
wire v$SEL5_15_out0;
wire v$SEL6_101_out0;
wire v$SEL6_132_out0;
wire v$SEL7_182_out0;
wire v$SEL7_94_out0;
wire v$SEL8_21_out0;
wire v$SEL9_35_out0;
wire v$SERIESCONNECT_193_out0;
wire v$SERIESCONNECT_289_out0;
wire v$_127_out1;

always @(posedge clk) v$REG1_103_out0 <= v$_51_out0;
always @(posedge clk) v$REG2_315_out0 <= v$INPUT_183_out0;
assign v$C19_330_out0 = 5'h9;
assign v$C3_328_out0 = 4'h1;
assign v$C13_326_out0 = 5'h1;
assign v$C21_324_out0 = 5'hb;
assign v$C6_298_out0 = 4'h4;
assign v$C5_284_out0 = 4'h3;
assign v$C2_283_out0 = 4'h0;
assign v$C1_276_out0 = 5'h2;
assign v$C30_274_out0 = 5'h14;
assign v$C11_263_out0 = 5'h3;
assign v$C18_250_out0 = 5'h11;
assign v$C10_239_out0 = 5'h0;
assign v$C31_229_out0 = 5'h13;
assign v$C11_208_out0 = 4'h9;
assign v$C4_203_out0 = 5'h8;
assign v$C8_189_out0 = 5'h7;
assign v$C9_171_out0 = 4'h7;
assign v$C14_168_out0 = 4'hc;
assign v$C8_161_out0 = 4'h6;
assign v$C12_146_out0 = 4'ha;
assign v$C1_145_out0 = 4'h0;
assign v$C15_135_out0 = 5'hd;
assign v$C10_125_out0 = 4'h8;
assign v$C7_123_out0 = 4'h5;
assign v$C20_95_out0 = 5'hc;
assign v$C3_93_out0 = 5'h5;
assign v$C12_92_out0 = 5'h4;
assign v$C13_90_out0 = 4'hb;
assign v$C17_75_out0 = 5'h10;
assign v$C4_68_out0 = 4'h2;
assign v$C28_67_out0 = 5'h12;
assign v$C14_43_out0 = 5'hf;
assign v$C16_27_out0 = 5'he;
assign v$C22_25_out0 = 5'ha;
assign v$C6_4_out0 = 5'h6;
assign v$_127_out0 = v$REG2_315_out0[20:0];
assign v$_127_out1 = v$REG2_315_out0[21:1];
assign v$OUTPUT_316_out0 = v$REG1_103_out0;
assign v$SEL8_21_out0 = v$OUTPUT_316_out0[8:8];
assign v$SEL9_35_out0 = v$OUTPUT_316_out0[0:0];
assign v$SEL16_79_out0 = v$OUTPUT_316_out0[15:15];
assign v$SEL22_88_out0 = v$OUTPUT_316_out0[14:14];
assign v$SEL5_124_out0 = v$OUTPUT_316_out0[2:2];
assign v$SEL6_132_out0 = v$OUTPUT_316_out0[12:12];
assign v$SEL1_151_out0 = v$OUTPUT_316_out0[5:5];
assign v$SEL2_154_out0 = v$OUTPUT_316_out0[3:3];
assign v$_157_out0 = v$_127_out0[7:0];
assign v$_157_out1 = v$_127_out0[20:13];
assign v$SEL11_158_out0 = v$OUTPUT_316_out0[10:10];
assign v$SEL7_182_out0 = v$OUTPUT_316_out0[11:11];
assign v$SEL26_197_out0 = v$OUTPUT_316_out0[19:19];
assign v$SEL19_202_out0 = v$OUTPUT_316_out0[16:16];
assign v$SEL10_215_out0 = v$OUTPUT_316_out0[1:1];
assign v$SEL18_221_out0 = v$OUTPUT_316_out0[18:18];
assign v$SEL12_249_out0 = v$OUTPUT_316_out0[9:9];
assign v$SEL13_252_out0 = v$OUTPUT_316_out0[4:4];
assign v$SEL25_269_out0 = v$OUTPUT_316_out0[20:20];
assign v$SEL3_295_out0 = v$OUTPUT_316_out0[7:7];
assign v$SEL24_299_out0 = v$OUTPUT_316_out0[17:17];
assign v$MSB_303_out0 = v$_127_out1;
assign v$SEL15_307_out0 = v$OUTPUT_316_out0[13:13];
assign v$SEL4_317_out0 = v$OUTPUT_316_out0[6:6];
assign v$4_5_out0 = v$SEL13_252_out0;
assign v$18_8_out0 = v$SEL18_221_out0;
assign v$15_16_out0 = v$SEL16_79_out0;
assign v$17_24_out0 = v$SEL24_299_out0;
assign v$19_34_out0 = v$SEL26_197_out0;
assign v$6_44_out0 = v$SEL4_317_out0;
assign v$5_49_out0 = v$SEL1_151_out0;
assign v$3_62_out0 = v$SEL2_154_out0;
assign v$7_70_out0 = v$SEL3_295_out0;
assign v$13_80_out0 = v$SEL15_307_out0;
assign v$2_97_out0 = v$SEL5_124_out0;
assign v$0_108_out0 = v$SEL9_35_out0;
assign v$10_114_out0 = v$SEL11_158_out0;
assign v$16_116_out0 = v$SEL19_202_out0;
assign v$1_121_out0 = v$SEL10_215_out0;
assign v$14_136_out0 = v$SEL22_88_out0;
assign v$9_176_out0 = v$SEL12_249_out0;
assign v$8_185_out0 = v$SEL8_21_out0;
assign v$12_188_out0 = v$SEL6_132_out0;
assign v$INPUT_190_out0 = v$_157_out1;
assign v$INPUT_191_out0 = v$_157_out0;
assign v$20_244_out0 = v$SEL25_269_out0;
assign v$11_313_out0 = v$SEL7_182_out0;
assign v$SEL18_2_out0 = v$INPUT_190_out0[3:3];
assign v$SEL18_3_out0 = v$INPUT_191_out0[3:3];
assign v$SEL5_15_out0 = v$INPUT_190_out0[10:10];
assign v$SEL15_28_out0 = v$INPUT_190_out0[4:4];
assign v$SEL15_29_out0 = v$INPUT_191_out0[4:4];
assign v$SEL14_77_out0 = v$INPUT_190_out0[7:7];
assign v$SEL14_78_out0 = v$INPUT_191_out0[7:7];
assign v$SEL12_81_out0 = v$INPUT_190_out0[12:12];
assign v$SEL7_94_out0 = v$INPUT_190_out0[8:8];
assign v$SEL6_101_out0 = v$INPUT_190_out0[9:9];
assign v$SEL21_133_out0 = v$INPUT_190_out0[0:0];
assign v$SEL21_134_out0 = v$INPUT_191_out0[0:0];
assign v$SEL20_140_out0 = v$INPUT_190_out0[1:1];
assign v$SEL20_141_out0 = v$INPUT_191_out0[1:1];
assign v$SEL13_223_out0 = v$INPUT_190_out0[6:6];
assign v$SEL13_224_out0 = v$INPUT_191_out0[6:6];
assign v$SEL17_259_out0 = v$INPUT_190_out0[2:2];
assign v$SEL17_260_out0 = v$INPUT_191_out0[2:2];
assign v$SEL16_266_out0 = v$INPUT_190_out0[5:5];
assign v$SEL16_267_out0 = v$INPUT_191_out0[5:5];
assign v$SEL1_294_out0 = v$INPUT_190_out0[11:11];
assign v$MUX4_331_out0 = v$20_244_out0 ? v$C10_239_out0 : v$C10_239_out0;
assign v$G52_17_out0 = ! v$SEL15_28_out0;
assign v$G52_18_out0 = ! v$SEL15_29_out0;
assign v$G66_40_out0 = ! v$SEL21_133_out0;
assign v$G46_41_out0 = ! v$SEL13_223_out0;
assign v$G46_42_out0 = ! v$SEL13_224_out0;
assign v$G19_52_out0 = ! v$SEL5_15_out0;
assign v$G17_72_out0 = ! v$SEL1_294_out0;
assign v$G39_91_out0 = ! v$SEL12_81_out0;
assign v$G40_142_out0 = ! v$SEL7_94_out0;
assign v$G45_169_out0 = ! v$SEL14_77_out0;
assign v$G45_170_out0 = ! v$SEL14_78_out0;
assign v$G22_207_out0 = ! v$SEL6_101_out0;
assign v$G51_232_out0 = ! v$SEL16_266_out0;
assign v$G51_233_out0 = ! v$SEL16_267_out0;
assign v$G58_287_out0 = ! v$SEL17_259_out0;
assign v$G58_288_out0 = ! v$SEL17_260_out0;
assign v$G57_301_out0 = ! v$SEL18_2_out0;
assign v$G57_302_out0 = ! v$SEL18_3_out0;
assign v$MUX12_304_out0 = v$19_34_out0 ? v$C13_326_out0 : v$MUX4_331_out0;
assign v$G62_305_out0 = ! v$SEL20_140_out0;
assign v$G62_306_out0 = ! v$SEL20_141_out0;
assign v$12_325_out0 = v$SEL12_81_out0;
assign v$MUX13_57_out0 = v$12_325_out0 ? v$C2_283_out0 : v$C1_145_out0;
assign v$MUX13_113_out0 = v$18_8_out0 ? v$C1_276_out0 : v$MUX12_304_out0;
assign v$G18_130_out0 = v$G17_72_out0 && v$G39_91_out0;
assign v$G6_212_out0 = v$SEL1_294_out0 && v$G39_91_out0;
assign v$G20_19_out0 = v$SEL5_15_out0 && v$G18_130_out0;
assign v$G23_100_out0 = v$G19_52_out0 && v$G18_130_out0;
assign v$11_275_out0 = v$G6_212_out0;
assign v$MUX2_327_out0 = v$17_24_out0 ? v$C11_263_out0 : v$MUX13_113_out0;
assign v$10_39_out0 = v$G20_19_out0;
assign v$MUX7_48_out0 = v$16_116_out0 ? v$C12_92_out0 : v$MUX2_327_out0;
assign v$G26_54_out0 = v$G22_207_out0 && v$G23_100_out0;
assign v$G21_115_out0 = v$SEL6_101_out0 && v$G23_100_out0;
assign v$MUX9_222_out0 = v$11_275_out0 ? v$C3_328_out0 : v$MUX13_57_out0;
assign v$_319_out0 = { v$12_325_out0,v$11_275_out0 };
assign v$9_160_out0 = v$G21_115_out0;
assign v$G24_164_out0 = v$SEL7_94_out0 && v$G26_54_out0;
assign v$G42_165_out0 = v$G40_142_out0 && v$G26_54_out0;
assign v$MUX12_251_out0 = v$10_39_out0 ? v$C4_68_out0 : v$MUX9_222_out0;
assign v$MUX8_265_out0 = v$15_16_out0 ? v$C3_93_out0 : v$MUX7_48_out0;
assign v$MUX10_45_out0 = v$9_160_out0 ? v$C5_284_out0 : v$MUX12_251_out0;
assign v$_71_out0 = { v$10_39_out0,v$9_160_out0 };
assign v$G41_98_out0 = v$G45_169_out0 && v$G42_165_out0;
assign v$8_126_out0 = v$G24_164_out0;
assign v$G43_155_out0 = v$SEL14_77_out0 && v$G42_165_out0;
assign v$MUX11_314_out0 = v$14_136_out0 ? v$C6_4_out0 : v$MUX8_265_out0;
assign v$MUX11_122_out0 = v$8_126_out0 ? v$C6_298_out0 : v$MUX10_45_out0;
assign v$G48_166_out0 = v$G46_41_out0 && v$G41_98_out0;
assign v$G44_200_out0 = v$SEL13_223_out0 && v$G41_98_out0;
assign v$MUX6_204_out0 = v$13_80_out0 ? v$C8_189_out0 : v$MUX11_314_out0;
assign v$_234_out0 = { v$_319_out0,v$_71_out0 };
assign v$7_308_out0 = v$G43_155_out0;
assign v$MUX1_33_out0 = v$12_188_out0 ? v$C4_203_out0 : v$MUX6_204_out0;
assign v$_109_out0 = { v$8_126_out0,v$7_308_out0 };
assign v$MUX8_150_out0 = v$7_308_out0 ? v$C7_123_out0 : v$MUX11_122_out0;
assign v$G49_216_out0 = v$SEL16_266_out0 && v$G48_166_out0;
assign v$6_227_out0 = v$G44_200_out0;
assign v$G47_279_out0 = v$G51_232_out0 && v$G48_166_out0;
assign v$G50_13_out0 = v$SEL15_28_out0 && v$G47_279_out0;
assign v$G54_128_out0 = v$G52_17_out0 && v$G47_279_out0;
assign v$MUX6_194_out0 = v$6_227_out0 ? v$C8_161_out0 : v$MUX8_150_out0;
assign v$5_270_out0 = v$G49_216_out0;
assign v$MUX22_333_out0 = v$11_313_out0 ? v$C19_330_out0 : v$MUX1_33_out0;
assign v$4_84_out0 = v$G50_13_out0;
assign v$MUX5_110_out0 = v$5_270_out0 ? v$C9_171_out0 : v$MUX6_194_out0;
assign v$MUX19_137_out0 = v$10_114_out0 ? v$C22_25_out0 : v$MUX22_333_out0;
assign v$G53_143_out0 = v$G57_301_out0 && v$G54_128_out0;
assign v$G55_213_out0 = v$SEL18_2_out0 && v$G54_128_out0;
assign v$_296_out0 = { v$6_227_out0,v$5_270_out0 };
assign v$MUX7_38_out0 = v$4_84_out0 ? v$C10_125_out0 : v$MUX5_110_out0;
assign v$G56_174_out0 = v$SEL17_259_out0 && v$G53_143_out0;
assign v$_195_out0 = { v$_109_out0,v$_296_out0 };
assign v$MUX16_264_out0 = v$9_176_out0 ? v$C21_324_out0 : v$MUX19_137_out0;
assign v$3_291_out0 = v$G55_213_out0;
assign v$G60_334_out0 = v$G58_287_out0 && v$G53_143_out0;
assign v$_0_out0 = { v$4_84_out0,v$3_291_out0 };
assign v$MUX4_50_out0 = v$3_291_out0 ? v$C11_208_out0 : v$MUX7_38_out0;
assign v$G63_55_out0 = v$G62_305_out0 && v$G60_334_out0;
assign v$_149_out0 = { v$_234_out0,v$_195_out0 };
assign v$2_177_out0 = v$G56_174_out0;
assign v$MUX21_256_out0 = v$8_185_out0 ? v$C20_95_out0 : v$MUX16_264_out0;
assign v$G61_257_out0 = v$SEL20_140_out0 && v$G60_334_out0;
assign v$G65_7_out0 = v$G66_40_out0 && v$G63_55_out0;
assign v$MUX15_96_out0 = v$7_70_out0 ? v$C15_135_out0 : v$MUX21_256_out0;
assign v$G64_162_out0 = v$G63_55_out0 && v$SEL21_133_out0;
assign v$MUX3_184_out0 = v$2_177_out0 ? v$C12_146_out0 : v$MUX4_50_out0;
assign v$1_219_out0 = v$G61_257_out0;
assign v$_22_out0 = { v$2_177_out0,v$1_219_out0 };
assign v$MUX2_69_out0 = v$1_219_out0 ? v$C13_90_out0 : v$MUX3_184_out0;
assign v$0_277_out0 = v$G64_162_out0;
assign v$SERIESCONNECT_289_out0 = v$G65_7_out0;
assign v$MUX18_332_out0 = v$6_44_out0 ? v$C16_27_out0 : v$MUX15_96_out0;
assign v$_30_out0 = { v$0_277_out0,v$1_219_out0 };
assign v$_65_out0 = { v$_0_out0,v$_22_out0 };
assign v$MUX1_179_out0 = v$0_277_out0 ? v$C14_168_out0 : v$MUX2_69_out0;
assign v$SERIESCONNECT_193_out0 = v$SERIESCONNECT_289_out0;
assign v$MUX20_268_out0 = v$5_49_out0 ? v$C14_43_out0 : v$MUX18_332_out0;
assign v$SHIFTNUMBER_20_out0 = v$MUX1_179_out0;
assign v$_82_out0 = { v$_30_out0,v$2_177_out0 };
assign v$G41_99_out0 = v$G45_170_out0 && v$SERIESCONNECT_193_out0;
assign v$G43_156_out0 = v$SEL14_78_out0 && v$SERIESCONNECT_193_out0;
assign v$MUX17_209_out0 = v$4_5_out0 ? v$C17_75_out0 : v$MUX20_268_out0;
assign v$_235_out0 = { v$_65_out0,v$0_277_out0 };
assign v$_152_out0 = { v$_149_out0,v$_235_out0 };
assign v$NOTUSE_159_out0 = v$SHIFTNUMBER_20_out0;
assign v$G48_167_out0 = v$G46_42_out0 && v$G41_99_out0;
assign v$MUX14_198_out0 = v$3_62_out0 ? v$C18_250_out0 : v$MUX17_209_out0;
assign v$G44_201_out0 = v$SEL13_224_out0 && v$G41_99_out0;
assign v$_237_out0 = { v$_82_out0,v$3_291_out0 };
assign v$7_309_out0 = v$G43_156_out0;
assign v$MUX31_104_out0 = v$2_97_out0 ? v$C28_67_out0 : v$MUX14_198_out0;
assign v$G49_217_out0 = v$SEL16_267_out0 && v$G48_167_out0;
assign v$6_228_out0 = v$G44_201_out0;
assign v$G47_280_out0 = v$G51_233_out0 && v$G48_167_out0;
assign v$_281_out0 = { v$_237_out0,v$4_84_out0 };
assign v$OUTPUTSHIFT_320_out0 = v$_152_out0;
assign v$G50_14_out0 = v$SEL15_29_out0 && v$G47_280_out0;
assign v$MUX28_53_out0 = v$1_121_out0 ? v$C31_229_out0 : v$MUX31_104_out0;
assign v$_86_out0 = { v$_281_out0,v$5_270_out0 };
assign v$NOTUSE1_102_out0 = v$OUTPUTSHIFT_320_out0;
assign v$G54_129_out0 = v$G52_18_out0 && v$G47_280_out0;
assign v$5_271_out0 = v$G49_217_out0;
assign v$_9_out0 = { v$_86_out0,v$6_227_out0 };
assign v$4_85_out0 = v$G50_14_out0;
assign v$G53_144_out0 = v$G57_302_out0 && v$G54_129_out0;
assign v$G55_214_out0 = v$SEL18_3_out0 && v$G54_129_out0;
assign v$_297_out0 = { v$6_228_out0,v$5_271_out0 };
assign v$MUX25_322_out0 = v$0_108_out0 ? v$C30_274_out0 : v$MUX28_53_out0;
assign v$G56_175_out0 = v$SEL17_260_out0 && v$G53_144_out0;
assign v$SHIFTNUMBER_186_out0 = v$MUX25_322_out0;
assign v$_196_out0 = { v$7_309_out0,v$_297_out0 };
assign v$_210_out0 = { v$_9_out0,v$7_308_out0 };
assign v$3_292_out0 = v$G55_214_out0;
assign v$G60_335_out0 = v$G58_288_out0 && v$G53_144_out0;
assign v$_1_out0 = { v$4_85_out0,v$3_292_out0 };
assign v$_6_out0 = { v$_210_out0,v$8_126_out0 };
assign v$G63_56_out0 = v$G62_306_out0 && v$G60_335_out0;
assign v$2_178_out0 = v$G56_175_out0;
assign v$G61_258_out0 = v$SEL20_141_out0 && v$G60_335_out0;
assign v$_89_out0 = { v$_6_out0,v$9_160_out0 };
assign v$G64_163_out0 = v$G63_56_out0 && v$SEL21_134_out0;
assign v$1_220_out0 = v$G61_258_out0;
assign v$_23_out0 = { v$2_178_out0,v$1_220_out0 };
assign v$_64_out0 = { v$_89_out0,v$10_39_out0 };
assign v$0_278_out0 = v$G64_163_out0;
assign v$_31_out0 = { v$0_278_out0,v$1_220_out0 };
assign v$_66_out0 = { v$_1_out0,v$_23_out0 };
assign v$_329_out0 = { v$_64_out0,v$11_275_out0 };
assign v$_47_out0 = { v$_329_out0,v$12_325_out0 };
assign v$_83_out0 = { v$_31_out0,v$2_178_out0 };
assign v$_236_out0 = { v$_66_out0,v$0_278_out0 };
assign v$OUTPUT_117_out0 = v$_47_out0;
assign v$_153_out0 = { v$_196_out0,v$_236_out0 };
assign v$_238_out0 = { v$_83_out0,v$3_292_out0 };
assign v$_282_out0 = { v$_238_out0,v$4_85_out0 };
assign v$OUTPUTSHIFT_321_out0 = v$_153_out0;
assign v$_87_out0 = { v$_282_out0,v$5_271_out0 };
assign v$NOTUSE2_241_out0 = v$OUTPUTSHIFT_321_out0;
assign v$_10_out0 = { v$_87_out0,v$6_228_out0 };
assign v$_211_out0 = { v$_10_out0,v$7_309_out0 };
assign v$OUTPUT_118_out0 = v$_211_out0;
assign v$_51_out0 = { v$OUTPUT_118_out0,v$OUTPUT_117_out0 };


endmodule
