

    module v$RAM3_1304(q, a, d, we, clk);
    output reg [15:0] q;
    input [15:0] d;
    input [11:0] a;
    input we, clk;
    reg [15:0] ram [4095:0];
     always @(posedge clk) begin
         if (we)
             ram[a] <= d;
         q <= ram[a];
     end

    integer i;
    initial
    begin
        for (i=0; i < 4096; i=i+1)
        begin
            ram[i] = 0;
        end

        ram[0] = 0;
ram[1792] = 15360;
ram[1793] = 12629;
ram[1794] = 0;
ram[1795] = 7236;
ram[1797] = 2688;
ram[1798] = 0;
    end
    endmodule

    

    module v$ROM3_3844(q, a, clk);
    output reg [15:0] q;
    input clk;
    input [11:0] a;
    reg [15:0] rom [4095:0];
    always @(posedge clk) q <= rom[a];
    integer i;
    initial
    begin
        for (i=0; i < 4096; i=i+1)
        begin
            rom[i] = 0;
        end
    
        rom[0] = 49799;
rom[1] = 50825;
rom[2] = 2884;
rom[3] = 3584;
rom[4] = 3265;
rom[5] = 2253;
rom[6] = 2253;
rom[7] = 2253;
rom[8] = 3793;
rom[9] = 3524;
rom[10] = 4036;
rom[11] = 3265;
rom[12] = 2253;
rom[13] = 2253;
rom[14] = 2253;
rom[15] = 2253;
rom[16] = 2253;
rom[17] = 3793;
rom[18] = 3524;
rom[19] = 4036;
rom[20] = 3265;
rom[21] = 2253;
rom[22] = 2253;
rom[23] = 2253;
rom[24] = 2253;
rom[25] = 2253;
rom[26] = 2253;
rom[27] = 2253;
rom[28] = 3793;
rom[29] = 3524;
rom[30] = 49799;
rom[31] = 2241;
rom[32] = 3016;
rom[33] = 2249;
rom[34] = 3016;
rom[35] = 2245;
rom[36] = 3016;
rom[37] = 2249;
rom[38] = 3792;
rom[39] = 3524;
rom[40] = 28672;
    end
    endmodule
     

    module v$ROM4_4954(q, a, clk);
    output reg [15:0] q;
    input clk;
    input [11:0] a;
    reg [15:0] rom [4095:0];
    always @(posedge clk) q <= rom[a];
    integer i;
    initial
    begin
        for (i=0; i < 4096; i=i+1)
        begin
            rom[i] = 0;
        end
    
        rom[0] = 49799;
rom[1] = 50825;
rom[2] = 2884;
rom[3] = 3584;
rom[4] = 3265;
rom[5] = 2253;
rom[6] = 2253;
rom[7] = 2253;
rom[8] = 3793;
rom[9] = 3524;
rom[10] = 4036;
rom[11] = 3265;
rom[12] = 2253;
rom[13] = 2253;
rom[14] = 2253;
rom[15] = 2253;
rom[16] = 2253;
rom[17] = 3793;
rom[18] = 3524;
rom[19] = 4036;
rom[20] = 3265;
rom[21] = 2253;
rom[22] = 2253;
rom[23] = 2253;
rom[24] = 2253;
rom[25] = 2253;
rom[26] = 2253;
rom[27] = 2253;
rom[28] = 3793;
rom[29] = 3524;
rom[30] = 49799;
rom[31] = 2241;
rom[32] = 3016;
rom[33] = 2249;
rom[34] = 3016;
rom[35] = 2245;
rom[36] = 3016;
rom[37] = 2249;
rom[38] = 3792;
rom[39] = 3524;
rom[40] = 28672;
    end
    endmodule
     
module main (
	clk,
	v$INTERRUPT2_976_out0,
	v$INTERRUPT1_3115_out0);
input clk;
input v$INTERRUPT1_3115_out0;
input v$INTERRUPT2_976_out0;
reg  [11:0] v$REG1_374_out0 = 12'h0;
reg  [11:0] v$REG1_375_out0 = 12'h0;
reg  [11:0] v$REG2_750_out0 = 12'h0;
reg  [11:0] v$REG2_751_out0 = 12'h0;
reg  [15:0] v$REG0_4539_out0 = 16'h0;
reg  [15:0] v$REG0_4540_out0 = 16'h0;
reg  [15:0] v$REG1_1106_out0 = 16'h0;
reg  [15:0] v$REG1_1399_out0 = 16'h0;
reg  [15:0] v$REG1_1400_out0 = 16'h0;
reg  [15:0] v$REG1_2682_out0 = 16'h0;
reg  [15:0] v$REG1_2683_out0 = 16'h0;
reg  [15:0] v$REG1_3272_out0 = 16'h0;
reg  [15:0] v$REG1_3273_out0 = 16'h0;
reg  [15:0] v$REG1_3653_out0 = 16'h0;
reg  [15:0] v$REG1_3654_out0 = 16'h0;
reg  [15:0] v$REG2_2762_out0 = 16'h0;
reg  [15:0] v$REG2_2763_out0 = 16'h0;
reg  [15:0] v$REG2_4872_out0 = 16'h0;
reg  [15:0] v$REG2_4873_out0 = 16'h0;
reg  [15:0] v$REG2_5309_out0 = 16'h0;
reg  [15:0] v$REG3_2164_out0 = 16'h0;
reg  [15:0] v$REG3_2165_out0 = 16'h0;
reg  [15:0] v$REG3_2962_out0 = 16'h0;
reg  [15:0] v$REG3_2963_out0 = 16'h0;
reg  [15:0] v$REG4_1772_out0 = 16'h0;
reg  [15:0] v$REG4_1773_out0 = 16'h0;
reg  [15:0] v$REG4_4843_out0 = 16'h0;
reg  [15:0] v$REG4_4844_out0 = 16'h0;
reg  [15:0] v$REG5_3036_out0 = 16'h0;
reg  [15:0] v$REG5_3037_out0 = 16'h0;
reg v$FF1_144_out0 = 1'b0;
reg v$FF1_145_out0 = 1'b0;
reg v$FF1_1575_out0 = 1'b0;
reg v$FF1_1576_out0 = 1'b0;
reg v$FF1_1618_out0 = 1'b0;
reg v$FF1_1619_out0 = 1'b0;
reg v$FF1_2042_out0 = 1'b0;
reg v$FF1_2043_out0 = 1'b0;
reg v$FF1_2233_out0 = 1'b0;
reg v$FF1_2975_out0 = 1'b0;
reg v$FF1_2976_out0 = 1'b0;
reg v$FF1_4133_out0 = 1'b0;
reg v$FF1_4134_out0 = 1'b0;
reg v$FF1_5073_out0 = 1'b0;
reg v$FF1_846_out0 = 1'b0;
reg v$FF2_1859_out0 = 1'b0;
reg v$FF2_2554_out0 = 1'b0;
reg v$FF2_2555_out0 = 1'b0;
reg v$FF2_3299_out0 = 1'b0;
reg v$FF2_3300_out0 = 1'b0;
reg v$FF2_3403_out0 = 1'b0;
reg v$FF2_4169_out0 = 1'b0;
reg v$FF2_4170_out0 = 1'b0;
reg v$FF2_4405_out0 = 1'b0;
reg v$FF2_4406_out0 = 1'b0;
reg v$FF3_4436_out0 = 1'b0;
reg v$FF3_4437_out0 = 1'b0;
reg v$FF4_3156_out0 = 1'b0;
reg v$FF4_3157_out0 = 1'b0;
reg v$FF4_89_out0 = 1'b0;
reg v$FF5_271_out0 = 1'b0;
reg v$REG2_1904_out0 = 1'b0;
reg v$REG2_1905_out0 = 1'b0;
reg v$REG3_574_out0 = 1'b0;
reg v$REG3_575_out0 = 1'b0;
wire  [10:0] v$A1_4358_out0;
wire  [10:0] v$A_1802_out0;
wire  [10:0] v$A_470_out0;
wire  [10:0] v$A_471_out0;
wire  [10:0] v$A_472_out0;
wire  [10:0] v$A_473_out0;
wire  [10:0] v$A_474_out0;
wire  [10:0] v$A_475_out0;
wire  [10:0] v$A_476_out0;
wire  [10:0] v$A_477_out0;
wire  [10:0] v$A_478_out0;
wire  [10:0] v$A_479_out0;
wire  [10:0] v$A_480_out0;
wire  [10:0] v$B0_4321_out0;
wire  [10:0] v$B0_90_out0;
wire  [10:0] v$B_951_out0;
wire  [10:0] v$C11_1736_out0;
wire  [10:0] v$C11_4416_out0;
wire  [10:0] v$C11_671_out0;
wire  [10:0] v$C1_1146_out0;
wire  [10:0] v$C1_1147_out0;
wire  [10:0] v$C1_1312_out0;
wire  [10:0] v$F1_4615_out0;
wire  [10:0] v$FRAC11A_154_out0;
wire  [10:0] v$FRAC11B_2912_out0;
wire  [10:0] v$FRACA_4929_out0;
wire  [10:0] v$FRACB_4130_out0;
wire  [10:0] v$MULTIPLICAND_5224_out0;
wire  [10:0] v$MULTIPLIER_1024_out0;
wire  [10:0] v$SIGNIFICANT_3533_out0;
wire  [10:0] v$TOBIGALU_1227_out0;
wire  [10:0] v$TOSHIFT_1120_out0;
wire  [10:0] v$X13_3686_out0;
wire  [10:0] v$X16_4534_out0;
wire  [10:0] v$X1_381_out0;
wire  [10:0] v$X1_382_out0;
wire  [10:0] v$X1_383_out0;
wire  [10:0] v$X1_384_out0;
wire  [10:0] v$X1_385_out0;
wire  [10:0] v$X1_386_out0;
wire  [10:0] v$X1_387_out0;
wire  [10:0] v$X1_388_out0;
wire  [10:0] v$X1_389_out0;
wire  [10:0] v$X1_390_out0;
wire  [10:0] v$X1_391_out0;
wire  [10:0] v$XOR2_4394_out0;
wire  [10:0] v$X_3_out0;
wire  [10:0] v$_1145_out0;
wire  [10:0] v$_1188_out0;
wire  [10:0] v$_1189_out0;
wire  [10:0] v$_1190_out0;
wire  [10:0] v$_1191_out0;
wire  [10:0] v$_1192_out0;
wire  [10:0] v$_1193_out0;
wire  [10:0] v$_1194_out0;
wire  [10:0] v$_1195_out0;
wire  [10:0] v$_1196_out0;
wire  [10:0] v$_1197_out0;
wire  [10:0] v$_1198_out0;
wire  [10:0] v$_1361_out1;
wire  [10:0] v$_1786_out0;
wire  [10:0] v$_196_out0;
wire  [10:0] v$_2070_out0;
wire  [10:0] v$_2401_out0;
wire  [10:0] v$_2687_out1;
wire  [10:0] v$_2944_out0;
wire  [10:0] v$_2993_out1;
wire  [10:0] v$_2994_out1;
wire  [10:0] v$_3051_out0;
wire  [10:0] v$_3067_out0;
wire  [10:0] v$_3067_out1;
wire  [10:0] v$_3580_out0;
wire  [10:0] v$_3710_out0;
wire  [10:0] v$_3831_out0;
wire  [10:0] v$_4536_out0;
wire  [10:0] v$_4748_out1;
wire  [10:0] v$_4940_out0;
wire  [10:0] v$_5099_out1;
wire  [10:0] v$_5100_out1;
wire  [10:0] v$_5251_out0;
wire  [10:0] v$_5259_out1;
wire  [10:0] v$_811_out0;
wire  [10:0] v$_933_out0;
wire  [10:0] v$_934_out0;
wire  [11:0] v$A1_2902_out0;
wire  [11:0] v$A1_2903_out0;
wire  [11:0] v$ADDRESS_1313_out0;
wire  [11:0] v$ADDRESS_2096_out0;
wire  [11:0] v$ADDRESS_4829_out0;
wire  [11:0] v$ADDRESS_4_out0;
wire  [11:0] v$B1_2488_out0;
wire  [11:0] v$B1_4597_out0;
wire  [11:0] v$C12_1162_out0;
wire  [11:0] v$C13_325_out0;
wire  [11:0] v$C1_1742_out0;
wire  [11:0] v$C1_1743_out0;
wire  [11:0] v$C1_2031_out0;
wire  [11:0] v$C1_2032_out0;
wire  [11:0] v$C4_3093_out0;
wire  [11:0] v$C4_3094_out0;
wire  [11:0] v$DATAADDRESS_2471_out0;
wire  [11:0] v$DATAADDRESS_2472_out0;
wire  [11:0] v$DMADDRESS_1885_out0;
wire  [11:0] v$IR110_4921_out0;
wire  [11:0] v$IR110_4922_out0;
wire  [11:0] v$IR12_3283_out0;
wire  [11:0] v$IR12_3284_out0;
wire  [11:0] v$LARGEREXP_3147_out0;
wire  [11:0] v$MUX1_3553_out0;
wire  [11:0] v$MUX1_3966_out0;
wire  [11:0] v$MUX1_3967_out0;
wire  [11:0] v$MUX2_1094_out0;
wire  [11:0] v$MUX2_769_out0;
wire  [11:0] v$MUX2_770_out0;
wire  [11:0] v$MUX4_2920_out0;
wire  [11:0] v$MUX4_788_out0;
wire  [11:0] v$MUX4_789_out0;
wire  [11:0] v$MUX5_2882_out0;
wire  [11:0] v$MUX5_2883_out0;
wire  [11:0] v$MUX5_3262_out0;
wire  [11:0] v$MUX6_3430_out0;
wire  [11:0] v$MUX6_3431_out0;
wire  [11:0] v$MUX7_4351_out0;
wire  [11:0] v$MUX7_4352_out0;
wire  [11:0] v$N_5020_out0;
wire  [11:0] v$N_5021_out0;
wire  [11:0] v$PC1_987_out0;
wire  [11:0] v$PC1_988_out0;
wire  [11:0] v$PC_4346_out0;
wire  [11:0] v$PC_4347_out0;
wire  [11:0] v$PROGRAMADDRESS_4514_out0;
wire  [11:0] v$PROGRAMADDRESS_4515_out0;
wire  [11:0] v$RAMADDRMUX_1479_out0;
wire  [11:0] v$RAMADDRMUX_1480_out0;
wire  [11:0] v$RAMADDRMUX_3785_out0;
wire  [11:0] v$RAMADDRMUX_3786_out0;
wire  [11:0] v$RAMADDRMUX_5262_out0;
wire  [11:0] v$RAMADDRMUX_5263_out0;
wire  [11:0] v$RAMADDRMUX_613_out0;
wire  [11:0] v$RAMADDRMUX_614_out0;
wire  [11:0] v$SMALLEREXP_3133_out0;
wire  [11:0] v$STOREDPC_3150_out0;
wire  [11:0] v$STOREDPC_3151_out0;
wire  [11:0] v$STOREDPC_5240_out0;
wire  [11:0] v$STOREDPC_5241_out0;
wire  [11:0] v$X16_4303_out0;
wire  [11:0] v$_1016_out1;
wire  [11:0] v$_1236_out1;
wire  [11:0] v$_1701_out1;
wire  [11:0] v$_1702_out1;
wire  [11:0] v$_1811_out0;
wire  [11:0] v$_1812_out1;
wire  [11:0] v$_1871_out1;
wire  [11:0] v$_2069_out0;
wire  [11:0] v$_2309_out0;
wire  [11:0] v$_2401_out1;
wire  [11:0] v$_2428_out1;
wire  [11:0] v$_2639_out1;
wire  [11:0] v$_2787_out1;
wire  [11:0] v$_2788_out1;
wire  [11:0] v$_3125_out1;
wire  [11:0] v$_3126_out1;
wire  [11:0] v$_3127_out1;
wire  [11:0] v$_3346_out0;
wire  [11:0] v$_3347_out0;
wire  [11:0] v$_3366_out1;
wire  [11:0] v$_3422_out0;
wire  [11:0] v$_3423_out0;
wire  [11:0] v$_3536_out0;
wire  [11:0] v$_3549_out0;
wire  [11:0] v$_3549_out1;
wire  [11:0] v$_3667_out1;
wire  [11:0] v$_3807_out1;
wire  [11:0] v$_3936_out0;
wire  [11:0] v$_4504_out0;
wire  [11:0] v$_4505_out0;
wire  [11:0] v$_4578_out1;
wire  [11:0] v$_4870_out1;
wire  [11:0] v$_4930_out0;
wire  [11:0] v$_503_out0;
wire  [11:0] v$_5398_out0;
wire  [11:0] v$_5399_out0;
wire  [11:0] v$_691_out1;
wire  [11:0] v$_861_out1;
wire  [12:0] v$0_1136_out0;
wire  [12:0] v$10_4736_out0;
wire  [12:0] v$11_3593_out0;
wire  [12:0] v$12_499_out0;
wire  [12:0] v$13_273_out0;
wire  [12:0] v$1_2087_out0;
wire  [12:0] v$2_320_out0;
wire  [12:0] v$3_1416_out0;
wire  [12:0] v$4_989_out0;
wire  [12:0] v$5_428_out0;
wire  [12:0] v$6_3566_out0;
wire  [12:0] v$7_129_out0;
wire  [12:0] v$8_3965_out0;
wire  [12:0] v$9_3469_out0;
wire  [12:0] v$A1_3679_out0;
wire  [12:0] v$ADD2_4212_out0;
wire  [12:0] v$B2_1401_out0;
wire  [12:0] v$B2_1666_out0;
wire  [12:0] v$C13_1012_out0;
wire  [12:0] v$C18_2405_out0;
wire  [12:0] v$C1_4937_out0;
wire  [12:0] v$C21_4143_out0;
wire  [12:0] v$C25_3774_out0;
wire  [12:0] v$C2_743_out0;
wire  [12:0] v$INPUT_3065_out0;
wire  [12:0] v$INPUT_3071_out0;
wire  [12:0] v$INPUT_3073_out0;
wire  [12:0] v$IN_1445_out0;
wire  [12:0] v$L0_2414_out0;
wire  [12:0] v$L1_2240_out0;
wire  [12:0] v$MUX10_1481_out0;
wire  [12:0] v$MUX11_2798_out0;
wire  [12:0] v$MUX12_3802_out0;
wire  [12:0] v$MUX13_3550_out0;
wire  [12:0] v$MUX14_1305_out0;
wire  [12:0] v$MUX15_5166_out0;
wire  [12:0] v$MUX17_1753_out0;
wire  [12:0] v$MUX18_2657_out0;
wire  [12:0] v$MUX19_1397_out0;
wire  [12:0] v$MUX1_3727_out0;
wire  [12:0] v$MUX1_4000_out0;
wire  [12:0] v$MUX20_3019_out0;
wire  [12:0] v$MUX21_779_out0;
wire  [12:0] v$MUX2_1808_out0;
wire  [12:0] v$MUX2_4855_out0;
wire  [12:0] v$MUX3_3189_out0;
wire  [12:0] v$MUX4_3470_out0;
wire  [12:0] v$MUX5_3232_out0;
wire  [12:0] v$MUX6_5236_out0;
wire  [12:0] v$MUX7_3999_out0;
wire  [12:0] v$MUX8_2088_out0;
wire  [12:0] v$MUX9_4512_out0;
wire  [12:0] v$NOTUSE1_1564_out0;
wire  [12:0] v$OUTPUTSHIFT_1089_out0;
wire  [12:0] v$OUTPUTSHIFT_5149_out0;
wire  [12:0] v$OUTPUTSHIFT_5151_out0;
wire  [12:0] v$OUTPUT_1819_out0;
wire  [12:0] v$OUTPUT_1821_out0;
wire  [12:0] v$OUTPUT_3581_out0;
wire  [12:0] v$OUTPUT_4621_out0;
wire  [12:0] v$SHIFTSIGNIFICANT_5041_out0;
wire  [12:0] v$SUM_5158_out0;
wire  [12:0] v$Toshift_5200_out0;
wire  [12:0] v$X21_241_out0;
wire  [12:0] v$XOR1_2651_out0;
wire  [12:0] v$X_1476_out0;
wire  [12:0] v$_1238_out1;
wire  [12:0] v$_1239_out1;
wire  [12:0] v$_1278_out0;
wire  [12:0] v$_1368_out0;
wire  [12:0] v$_1387_out1;
wire  [12:0] v$_1411_out0;
wire  [12:0] v$_1523_out0;
wire  [12:0] v$_1549_out0;
wire  [12:0] v$_164_out0;
wire  [12:0] v$_1770_out0;
wire  [12:0] v$_2027_out0;
wire  [12:0] v$_2196_out1;
wire  [12:0] v$_2197_out1;
wire  [12:0] v$_2235_out0;
wire  [12:0] v$_2423_out0;
wire  [12:0] v$_2425_out0;
wire  [12:0] v$_2501_out0;
wire  [12:0] v$_2516_out1;
wire  [12:0] v$_2637_out0;
wire  [12:0] v$_2750_out0;
wire  [12:0] v$_2755_out0;
wire  [12:0] v$_2837_out0;
wire  [12:0] v$_2939_out0;
wire  [12:0] v$_3000_out0;
wire  [12:0] v$_3003_out1;
wire  [12:0] v$_3050_out0;
wire  [12:0] v$_3560_out0;
wire  [12:0] v$_3860_out0;
wire  [12:0] v$_3901_out0;
wire  [12:0] v$_4008_out0;
wire  [12:0] v$_4638_out0;
wire  [12:0] v$_4730_out0;
wire  [12:0] v$_4828_out0;
wire  [12:0] v$_5254_out0;
wire  [12:0] v$_600_out0;
wire  [12:0] v$_601_out0;
wire  [12:0] v$_607_out0;
wire  [12:0] v$_771_out0;
wire  [13:0] v$B3_3095_out0;
wire  [13:0] v$B3_692_out0;
wire  [13:0] v$C28_4909_out0;
wire  [13:0] v$M0_573_out0;
wire  [13:0] v$X24_2269_out0;
wire  [13:0] v$_1080_out0;
wire  [13:0] v$_1081_out0;
wire  [13:0] v$_11_out1;
wire  [13:0] v$_12_out1;
wire  [13:0] v$_1728_out1;
wire  [13:0] v$_1729_out1;
wire  [13:0] v$_222_out0;
wire  [13:0] v$_3090_out0;
wire  [13:0] v$_3442_out0;
wire  [13:0] v$_3554_out0;
wire  [13:0] v$_3556_out1;
wire  [13:0] v$_3792_out0;
wire  [13:0] v$_4072_out0;
wire  [13:0] v$_4408_out1;
wire  [13:0] v$_4409_out1;
wire  [13:0] v$_5179_out0;
wire  [13:0] v$_747_out1;
wire  [14:0] v$A1_794_out0;
wire  [14:0] v$B4_380_out0;
wire  [14:0] v$B4_4037_out0;
wire  [14:0] v$C24_4122_out0;
wire  [14:0] v$SEL52_1439_out0;
wire  [14:0] v$SEL53_3630_out0;
wire  [14:0] v$X22_626_out0;
wire  [14:0] v$_1688_out1;
wire  [14:0] v$_1900_out0;
wire  [14:0] v$_2284_out0;
wire  [14:0] v$_2285_out0;
wire  [14:0] v$_256_out1;
wire  [14:0] v$_257_out1;
wire  [14:0] v$_2774_out0;
wire  [14:0] v$_3020_out0;
wire  [14:0] v$_328_out0;
wire  [14:0] v$_3534_out0;
wire  [14:0] v$_3535_out0;
wire  [14:0] v$_3772_out1;
wire  [14:0] v$_3773_out1;
wire  [14:0] v$_3784_out0;
wire  [14:0] v$_4095_out1;
wire  [14:0] v$_4372_out0;
wire  [14:0] v$_4683_out0;
wire  [14:0] v$_4906_out1;
wire  [14:0] v$_4907_out1;
wire  [14:0] v$_517_out0;
wire  [14:0] v$_880_out1;
wire  [14:0] v$_881_out1;
wire  [15:0] v$1TO4_3665_out0;
wire  [15:0] v$1TO4_3666_out0;
wire  [15:0] v$A1_1123_out0;
wire  [15:0] v$A1_1124_out0;
wire  [15:0] v$A1_331_out0;
wire  [15:0] v$A1_332_out0;
wire  [15:0] v$ALUOUT_1496_out0;
wire  [15:0] v$ALUOUT_1497_out0;
wire  [15:0] v$ALUOUT_1768_out0;
wire  [15:0] v$ALUOUT_1769_out0;
wire  [15:0] v$ALUOUT_3587_out0;
wire  [15:0] v$ALUOUT_3588_out0;
wire  [15:0] v$ALUOUT_3789_out0;
wire  [15:0] v$ALUOUT_3790_out0;
wire  [15:0] v$ALUOUT_5256_out0;
wire  [15:0] v$ALUOUT_5257_out0;
wire  [15:0] v$ALUOUT_545_out0;
wire  [15:0] v$ALUOUT_546_out0;
wire  [15:0] v$ANDOUT_3462_out0;
wire  [15:0] v$ANDOUT_3463_out0;
wire  [15:0] v$ASR_232_out0;
wire  [15:0] v$ASR_233_out0;
wire  [15:0] v$ASR_2947_out0;
wire  [15:0] v$ASR_2948_out0;
wire  [15:0] v$ASR_628_out0;
wire  [15:0] v$ASR_629_out0;
wire  [15:0] v$ASR_834_out0;
wire  [15:0] v$ASR_835_out0;
wire  [15:0] v$A_2331_out0;
wire  [15:0] v$A_4810_out0;
wire  [15:0] v$A_4811_out0;
wire  [15:0] v$A_5334_out0;
wire  [15:0] v$A_602_out0;
wire  [15:0] v$A_749_out0;
wire  [15:0] v$B5_2508_out0;
wire  [15:0] v$B5_3091_out0;
wire  [15:0] v$B_2005_out0;
wire  [15:0] v$B_3539_out0;
wire  [15:0] v$B_4103_out0;
wire  [15:0] v$B_4104_out0;
wire  [15:0] v$B_5057_out0;
wire  [15:0] v$B_5337_out0;
wire  [15:0] v$C1_864_out0;
wire  [15:0] v$C1_865_out0;
wire  [15:0] v$C2_5403_out0;
wire  [15:0] v$C2_5404_out0;
wire  [15:0] v$C30_3636_out0;
wire  [15:0] v$C3_1545_out0;
wire  [15:0] v$C3_1546_out0;
wire  [15:0] v$C4_395_out0;
wire  [15:0] v$C4_396_out0;
wire  [15:0] v$DATA_968_out0;
wire  [15:0] v$DIN3_3861_out0;
wire  [15:0] v$DIN3_3862_out0;
wire  [15:0] v$DM1_492_out0;
wire  [15:0] v$DM1_492_out1;
wire  [15:0] v$DM2_3561_out0;
wire  [15:0] v$DM2_3561_out1;
wire  [15:0] v$DMDATA_4516_out0;
wire  [15:0] v$DMDATA_5169_out0;
wire  [15:0] v$DOUT1_873_out0;
wire  [15:0] v$DOUT1_874_out0;
wire  [15:0] v$DOUT2_1013_out0;
wire  [15:0] v$DOUT2_1014_out0;
wire  [15:0] v$EA_2692_out0;
wire  [15:0] v$EA_2693_out0;
wire  [15:0] v$FPOUT_4289_out0;
wire  [15:0] v$FPOUT_4479_out0;
wire  [15:0] v$FPOUT_4831_out0;
wire  [15:0] v$IN_1026_out0;
wire  [15:0] v$IN_1027_out0;
wire  [15:0] v$IN_1798_out0;
wire  [15:0] v$IN_1799_out0;
wire  [15:0] v$IN_2394_out0;
wire  [15:0] v$IN_2395_out0;
wire  [15:0] v$IN_2403_out0;
wire  [15:0] v$IN_2404_out0;
wire  [15:0] v$IN_2966_out0;
wire  [15:0] v$IN_2967_out0;
wire  [15:0] v$IN_3131_out0;
wire  [15:0] v$IN_3132_out0;
wire  [15:0] v$IN_353_out0;
wire  [15:0] v$IN_354_out0;
wire  [15:0] v$IN_4526_out0;
wire  [15:0] v$IN_4527_out0;
wire  [15:0] v$IN_4576_out0;
wire  [15:0] v$IN_4577_out0;
wire  [15:0] v$IN_4895_out0;
wire  [15:0] v$IN_4896_out0;
wire  [15:0] v$IN_4914_out0;
wire  [15:0] v$IN_4915_out0;
wire  [15:0] v$IR16_5206_out0;
wire  [15:0] v$IR16_5207_out0;
wire  [15:0] v$IR_2357_out0;
wire  [15:0] v$IR_2358_out0;
wire  [15:0] v$IR_2617_out0;
wire  [15:0] v$IR_2618_out0;
wire  [15:0] v$IR_269_out0;
wire  [15:0] v$IR_270_out0;
wire  [15:0] v$IR_3909_out0;
wire  [15:0] v$IR_3910_out0;
wire  [15:0] v$IR_837_out0;
wire  [15:0] v$IR_838_out0;
wire  [15:0] v$L2_3025_out0;
wire  [15:0] v$L3_5181_out0;
wire  [15:0] v$LSL_1395_out0;
wire  [15:0] v$LSL_1396_out0;
wire  [15:0] v$LSL_2051_out0;
wire  [15:0] v$LSL_2052_out0;
wire  [15:0] v$LSL_3834_out0;
wire  [15:0] v$LSL_3835_out0;
wire  [15:0] v$LSL_5349_out0;
wire  [15:0] v$LSL_5350_out0;
wire  [15:0] v$LSR_2177_out0;
wire  [15:0] v$LSR_2178_out0;
wire  [15:0] v$LSR_2641_out0;
wire  [15:0] v$LSR_2642_out0;
wire  [15:0] v$LSR_3076_out0;
wire  [15:0] v$LSR_3077_out0;
wire  [15:0] v$LSR_4948_out0;
wire  [15:0] v$LSR_4949_out0;
wire  [15:0] v$M1_973_out0;
wire  [15:0] v$MSL_591_out0;
wire  [15:0] v$MSL_592_out0;
wire  [15:0] v$MSR_2502_out0;
wire  [15:0] v$MSR_2503_out0;
wire  [15:0] v$MUX10_2171_out0;
wire  [15:0] v$MUX10_2172_out0;
wire  [15:0] v$MUX11_1403_out0;
wire  [15:0] v$MUX11_1404_out0;
wire  [15:0] v$MUX12_152_out0;
wire  [15:0] v$MUX12_153_out0;
wire  [15:0] v$MUX13_4054_out0;
wire  [15:0] v$MUX13_4055_out0;
wire  [15:0] v$MUX14_1674_out0;
wire  [15:0] v$MUX14_1675_out0;
wire  [15:0] v$MUX1_1219_out0;
wire  [15:0] v$MUX1_1435_out0;
wire  [15:0] v$MUX1_1436_out0;
wire  [15:0] v$MUX1_1624_out0;
wire  [15:0] v$MUX1_1625_out0;
wire  [15:0] v$MUX1_2744_out0;
wire  [15:0] v$MUX1_2745_out0;
wire  [15:0] v$MUX1_3023_out0;
wire  [15:0] v$MUX1_3024_out0;
wire  [15:0] v$MUX1_3564_out0;
wire  [15:0] v$MUX1_3565_out0;
wire  [15:0] v$MUX1_3674_out0;
wire  [15:0] v$MUX1_3675_out0;
wire  [15:0] v$MUX1_3811_out0;
wire  [15:0] v$MUX1_3812_out0;
wire  [15:0] v$MUX1_3902_out0;
wire  [15:0] v$MUX1_3903_out0;
wire  [15:0] v$MUX1_3947_out0;
wire  [15:0] v$MUX1_4052_out0;
wire  [15:0] v$MUX1_4053_out0;
wire  [15:0] v$MUX1_4389_out0;
wire  [15:0] v$MUX1_4390_out0;
wire  [15:0] v$MUX1_4868_out0;
wire  [15:0] v$MUX1_4869_out0;
wire  [15:0] v$MUX1_5298_out0;
wire  [15:0] v$MUX1_5299_out0;
wire  [15:0] v$MUX2_2109_out0;
wire  [15:0] v$MUX2_2110_out0;
wire  [15:0] v$MUX2_2169_out0;
wire  [15:0] v$MUX2_2170_out0;
wire  [15:0] v$MUX2_2255_out0;
wire  [15:0] v$MUX2_2256_out0;
wire  [15:0] v$MUX2_2857_out0;
wire  [15:0] v$MUX2_2858_out0;
wire  [15:0] v$MUX2_3809_out0;
wire  [15:0] v$MUX2_3810_out0;
wire  [15:0] v$MUX2_4708_out0;
wire  [15:0] v$MUX2_4709_out0;
wire  [15:0] v$MUX2_5187_out0;
wire  [15:0] v$MUX2_792_out0;
wire  [15:0] v$MUX2_793_out0;
wire  [15:0] v$MUX3_2384_out0;
wire  [15:0] v$MUX3_2385_out0;
wire  [15:0] v$MUX3_3205_out0;
wire  [15:0] v$MUX3_3206_out0;
wire  [15:0] v$MUX3_3233_out0;
wire  [15:0] v$MUX3_3234_out0;
wire  [15:0] v$MUX3_3333_out0;
wire  [15:0] v$MUX3_3334_out0;
wire  [15:0] v$MUX3_366_out0;
wire  [15:0] v$MUX3_367_out0;
wire  [15:0] v$MUX3_462_out0;
wire  [15:0] v$MUX3_463_out0;
wire  [15:0] v$MUX3_4904_out0;
wire  [15:0] v$MUX3_4905_out0;
wire  [15:0] v$MUX3_5264_out0;
wire  [15:0] v$MUX3_5265_out0;
wire  [15:0] v$MUX3_5300_out0;
wire  [15:0] v$MUX4_1067_out0;
wire  [15:0] v$MUX4_1068_out0;
wire  [15:0] v$MUX4_1306_out0;
wire  [15:0] v$MUX4_1307_out0;
wire  [15:0] v$MUX4_1893_out0;
wire  [15:0] v$MUX4_1894_out0;
wire  [15:0] v$MUX4_276_out0;
wire  [15:0] v$MUX4_277_out0;
wire  [15:0] v$MUX4_407_out0;
wire  [15:0] v$MUX4_408_out0;
wire  [15:0] v$MUX4_413_out0;
wire  [15:0] v$MUX4_414_out0;
wire  [15:0] v$MUX4_5267_out0;
wire  [15:0] v$MUX4_5268_out0;
wire  [15:0] v$MUX4_936_out0;
wire  [15:0] v$MUX5_3080_out0;
wire  [15:0] v$MUX5_3081_out0;
wire  [15:0] v$MUX5_3743_out0;
wire  [15:0] v$MUX5_3744_out0;
wire  [15:0] v$MUX6_1469_out0;
wire  [15:0] v$MUX6_1470_out0;
wire  [15:0] v$MUX6_796_out0;
wire  [15:0] v$MUX6_797_out0;
wire  [15:0] v$MUX7_3001_out0;
wire  [15:0] v$MUX7_3002_out0;
wire  [15:0] v$MUX8_1725_out0;
wire  [15:0] v$MUX8_1726_out0;
wire  [15:0] v$MUX9_3795_out0;
wire  [15:0] v$MUX9_3796_out0;
wire  [15:0] v$OP1_1525_out0;
wire  [15:0] v$OP1_1526_out0;
wire  [15:0] v$OP1_4087_out0;
wire  [15:0] v$OP1_4088_out0;
wire  [15:0] v$OP2_2123_out0;
wire  [15:0] v$OP2_2124_out0;
wire  [15:0] v$OP2_2722_out0;
wire  [15:0] v$OP2_2723_out0;
wire  [15:0] v$OP2_2995_out0;
wire  [15:0] v$OP2_2996_out0;
wire  [15:0] v$OP2_4043_out0;
wire  [15:0] v$OP2_4044_out0;
wire  [15:0] v$OUT_1077_out0;
wire  [15:0] v$OUT_1078_out0;
wire  [15:0] v$OUT_1757_out0;
wire  [15:0] v$OUT_1758_out0;
wire  [15:0] v$OUT_3063_out0;
wire  [15:0] v$OUT_3064_out0;
wire  [15:0] v$OUT_4569_out0;
wire  [15:0] v$OUT_4570_out0;
wire  [15:0] v$OUT_5294_out0;
wire  [15:0] v$OUT_5295_out0;
wire  [15:0] v$PCORROM_3465_out0;
wire  [15:0] v$PCORROM_3466_out0;
wire  [15:0] v$R01_3542_out0;
wire  [15:0] v$R02_2546_out0;
wire  [15:0] v$R0S_1142_out0;
wire  [15:0] v$R0S_1143_out0;
wire  [15:0] v$R0S_1231_out0;
wire  [15:0] v$R0S_1232_out0;
wire  [15:0] v$R0TEST_2264_out0;
wire  [15:0] v$R0TEST_2265_out0;
wire  [15:0] v$R0TEST_5113_out0;
wire  [15:0] v$R0TEST_5114_out0;
wire  [15:0] v$R0_1056_out0;
wire  [15:0] v$R0_1057_out0;
wire  [15:0] v$R0_3873_out0;
wire  [15:0] v$R0_3874_out0;
wire  [15:0] v$R0_3907_out0;
wire  [15:0] v$R0_3908_out0;
wire  [15:0] v$R0_4215_out0;
wire  [15:0] v$R0_4216_out0;
wire  [15:0] v$R0_925_out0;
wire  [15:0] v$R0_926_out0;
wire  [15:0] v$R11_3434_out0;
wire  [15:0] v$R12_4500_out0;
wire  [15:0] v$R1S_279_out0;
wire  [15:0] v$R1S_280_out0;
wire  [15:0] v$R1S_4900_out0;
wire  [15:0] v$R1S_4901_out0;
wire  [15:0] v$R1TEST_2942_out0;
wire  [15:0] v$R1TEST_2943_out0;
wire  [15:0] v$R1TEST_4069_out0;
wire  [15:0] v$R1TEST_4070_out0;
wire  [15:0] v$R1_2934_out0;
wire  [15:0] v$R1_2935_out0;
wire  [15:0] v$R1_3682_out0;
wire  [15:0] v$R1_3683_out0;
wire  [15:0] v$R1_4116_out0;
wire  [15:0] v$R1_4117_out0;
wire  [15:0] v$R1_4338_out0;
wire  [15:0] v$R1_4339_out0;
wire  [15:0] v$R1_5052_out0;
wire  [15:0] v$R1_5053_out0;
wire  [15:0] v$R21_2715_out0;
wire  [15:0] v$R22_2273_out0;
wire  [15:0] v$R2S_1379_out0;
wire  [15:0] v$R2S_1380_out0;
wire  [15:0] v$R2S_3521_out0;
wire  [15:0] v$R2S_3522_out0;
wire  [15:0] v$R2TEST_1284_out0;
wire  [15:0] v$R2TEST_1285_out0;
wire  [15:0] v$R2TEST_4286_out0;
wire  [15:0] v$R2TEST_4287_out0;
wire  [15:0] v$R2_2167_out0;
wire  [15:0] v$R2_2168_out0;
wire  [15:0] v$R2_2904_out0;
wire  [15:0] v$R2_2905_out0;
wire  [15:0] v$R2_3009_out0;
wire  [15:0] v$R2_3010_out0;
wire  [15:0] v$R2_3953_out0;
wire  [15:0] v$R2_3954_out0;
wire  [15:0] v$R2_5037_out0;
wire  [15:0] v$R2_5038_out0;
wire  [15:0] v$R31_2229_out0;
wire  [15:0] v$R32_3176_out0;
wire  [15:0] v$R3S_4759_out0;
wire  [15:0] v$R3S_4760_out0;
wire  [15:0] v$R3S_4764_out0;
wire  [15:0] v$R3S_4765_out0;
wire  [15:0] v$R3TEST_2015_out0;
wire  [15:0] v$R3TEST_2016_out0;
wire  [15:0] v$R3TEST_5310_out0;
wire  [15:0] v$R3TEST_5311_out0;
wire  [15:0] v$R3_1883_out0;
wire  [15:0] v$R3_1884_out0;
wire  [15:0] v$R3_2053_out0;
wire  [15:0] v$R3_2054_out0;
wire  [15:0] v$R3_2227_out0;
wire  [15:0] v$R3_2228_out0;
wire  [15:0] v$R3_2875_out0;
wire  [15:0] v$R3_2876_out0;
wire  [15:0] v$R3_5058_out0;
wire  [15:0] v$R3_5059_out0;
wire  [15:0] v$RAM3_1304_out0;
wire  [15:0] v$RAMDOUT_2103_out0;
wire  [15:0] v$RAMDOUT_2104_out0;
wire  [15:0] v$RAMDOUT_2667_out0;
wire  [15:0] v$RAMDOUT_2668_out0;
wire  [15:0] v$RAMDOUT_2768_out0;
wire  [15:0] v$RAMDOUT_2769_out0;
wire  [15:0] v$RAMDOUT_2885_out0;
wire  [15:0] v$RAMDOUT_2886_out0;
wire  [15:0] v$RAMDOUT_4700_out0;
wire  [15:0] v$RAMDOUT_4701_out0;
wire  [15:0] v$RAMOUT_2337_out0;
wire  [15:0] v$RDOUT_1775_out0;
wire  [15:0] v$RDOUT_1776_out0;
wire  [15:0] v$RDOUT_289_out0;
wire  [15:0] v$RDOUT_290_out0;
wire  [15:0] v$RD_2135_out0;
wire  [15:0] v$RD_2136_out0;
wire  [15:0] v$READDATA1_2193_out0;
wire  [15:0] v$READDATA1_3559_out0;
wire  [15:0] v$READDATA2_2400_out0;
wire  [15:0] v$READDATA2_3664_out0;
wire  [15:0] v$REGDIN_1934_out0;
wire  [15:0] v$REGDIN_1935_out0;
wire  [15:0] v$REGDIN_3350_out0;
wire  [15:0] v$REGDIN_3351_out0;
wire  [15:0] v$RMN_3404_out0;
wire  [15:0] v$RMN_3405_out0;
wire  [15:0] v$RMN_844_out0;
wire  [15:0] v$RMN_845_out0;
wire  [15:0] v$RM_1148_out0;
wire  [15:0] v$RM_1149_out0;
wire  [15:0] v$RM_1744_out0;
wire  [15:0] v$RM_1745_out0;
wire  [15:0] v$RM_2274_out0;
wire  [15:0] v$RM_2275_out0;
wire  [15:0] v$RM_3021_out0;
wire  [15:0] v$RM_3022_out0;
wire  [15:0] v$RM_3453_out0;
wire  [15:0] v$RM_3454_out0;
wire  [15:0] v$RM_4530_out0;
wire  [15:0] v$RM_4531_out0;
wire  [15:0] v$RM_5033_out0;
wire  [15:0] v$RM_5034_out0;
wire  [15:0] v$ROM3_3844_out0;
wire  [15:0] v$ROM4_4954_out0;
wire  [15:0] v$ROR_1018_out0;
wire  [15:0] v$ROR_1019_out0;
wire  [15:0] v$ROR_1686_out0;
wire  [15:0] v$ROR_1687_out0;
wire  [15:0] v$ROR_2513_out0;
wire  [15:0] v$ROR_2514_out0;
wire  [15:0] v$ROR_2757_out0;
wire  [15:0] v$ROR_2758_out0;
wire  [15:0] v$SHIFTIN_2366_out0;
wire  [15:0] v$SHIFTIN_2367_out0;
wire  [15:0] v$SHIFTOUT_1795_out0;
wire  [15:0] v$SHIFTOUT_1796_out0;
wire  [15:0] v$WDATA_1785_out0;
wire  [15:0] v$WDATA_4407_out0;
wire  [15:0] v$WDATA_964_out0;
wire  [15:0] v$WDATA_965_out0;
wire  [15:0] v$WRITEDATA_1247_out0;
wire  [15:0] v$WRITEDATA_1248_out0;
wire  [15:0] v$WRITEDATA_1328_out0;
wire  [15:0] v$WRITEDATA_813_out0;
wire  [15:0] v$X27_3311_out0;
wire  [15:0] v$XOR1_1447_out0;
wire  [15:0] v$XOR1_1448_out0;
wire  [15:0] v$XOR1_2094_out0;
wire  [15:0] v$XOR1_2095_out0;
wire  [15:0] v$X_4521_out0;
wire  [15:0] v$X_4522_out0;
wire  [15:0] v$_1236_out0;
wire  [15:0] v$_1449_out0;
wire  [15:0] v$_1536_out0;
wire  [15:0] v$_1551_out0;
wire  [15:0] v$_1552_out0;
wire  [15:0] v$_1816_out0;
wire  [15:0] v$_1817_out0;
wire  [15:0] v$_19_out0;
wire  [15:0] v$_2089_out0;
wire  [15:0] v$_220_out0;
wire  [15:0] v$_221_out0;
wire  [15:0] v$_2440_out0;
wire  [15:0] v$_2484_out0;
wire  [15:0] v$_2485_out0;
wire  [15:0] v$_2578_out0;
wire  [15:0] v$_281_out0;
wire  [15:0] v$_282_out0;
wire  [15:0] v$_3045_out0;
wire  [15:0] v$_3046_out0;
wire  [15:0] v$_3061_out0;
wire  [15:0] v$_3062_out0;
wire  [15:0] v$_3101_out0;
wire  [15:0] v$_3102_out0;
wire  [15:0] v$_3415_out0;
wire  [15:0] v$_3416_out0;
wire  [15:0] v$_3447_out0;
wire  [15:0] v$_3448_out0;
wire  [15:0] v$_3641_out0;
wire  [15:0] v$_3642_out0;
wire  [15:0] v$_377_out0;
wire  [15:0] v$_378_out0;
wire  [15:0] v$_3799_out0;
wire  [15:0] v$_3800_out0;
wire  [15:0] v$_4151_out0;
wire  [15:0] v$_4152_out0;
wire  [15:0] v$_4153_out0;
wire  [15:0] v$_4154_out0;
wire  [15:0] v$_4564_out0;
wire  [15:0] v$_4691_out1;
wire  [15:0] v$_5152_out0;
wire  [15:0] v$_515_out0;
wire  [15:0] v$_5167_out1;
wire  [15:0] v$_516_out0;
wire  [15:0] v$_5287_out0;
wire  [15:0] v$_5288_out0;
wire  [15:0] v$_593_out0;
wire  [15:0] v$_594_out0;
wire  [15:0] v$_636_out0;
wire  [15:0] v$_637_out0;
wire  [15:0] v$_948_out0;
wire  [15:0] v$_949_out0;
wire  [15:0] v$_956_out0;
wire  [15:0] v$_957_out0;
wire  [15:0] v$fpmerge_5196_out0;
wire  [16:0] v$B6_2056_out0;
wire  [16:0] v$B6_262_out0;
wire  [16:0] v$C26_791_out0;
wire  [16:0] v$N0_1483_out0;
wire  [16:0] v$N0_1845_out0;
wire  [16:0] v$N0_3504_out0;
wire  [16:0] v$X18_2941_out0;
wire  [16:0] v$_1046_out1;
wire  [16:0] v$_3740_out0;
wire  [16:0] v$_3813_out0;
wire  [16:0] v$_4475_out1;
wire  [16:0] v$_4747_out0;
wire  [16:0] v$_4752_out0;
wire  [16:0] v$_5390_out0;
wire  [16:0] v$_735_out0;
wire  [17:0] v$B7_1140_out0;
wire  [17:0] v$B7_3060_out0;
wire  [17:0] v$C22_4676_out0;
wire  [17:0] v$X31_4020_out0;
wire  [17:0] v$_104_out0;
wire  [17:0] v$_3618_out0;
wire  [17:0] v$_365_out1;
wire  [17:0] v$_3677_out1;
wire  [17:0] v$_4579_out0;
wire  [18:0] v$B8_1901_out0;
wire  [18:0] v$B8_2200_out0;
wire  [18:0] v$C29_4076_out0;
wire  [18:0] v$L4_5246_out0;
wire  [18:0] v$L5_1655_out0;
wire  [18:0] v$M2_1829_out0;
wire  [18:0] v$N1_2746_out0;
wire  [18:0] v$N1_3180_out0;
wire  [18:0] v$N1_5023_out0;
wire  [18:0] v$X38_1004_out0;
wire  [18:0] v$_1240_out0;
wire  [18:0] v$_1371_out0;
wire  [18:0] v$_1716_out0;
wire  [18:0] v$_3525_out0;
wire  [18:0] v$_4532_out0;
wire  [18:0] v$_4862_out1;
wire  [18:0] v$_500_out0;
wire  [18:0] v$_8_out0;
wire  [18:0] v$_972_out1;
wire  [19:0] v$0_5061_out0;
wire  [19:0] v$B9_1681_out0;
wire  [19:0] v$B9_812_out0;
wire  [19:0] v$C25_3012_out0;
wire  [19:0] v$M3_3543_out0;
wire  [19:0] v$X20_2699_out0;
wire  [19:0] v$_1370_out0;
wire  [19:0] v$_1705_out0;
wire  [19:0] v$_2097_out1;
wire  [19:0] v$_2987_out0;
wire  [19:0] v$_3589_out0;
wire  [19:0] v$_4931_out1;
wire  [19:0] v$_950_out0;
wire  [1:0] v$2_3526_out0;
wire  [1:0] v$2_3527_out0;
wire  [1:0] v$3_31_out0;
wire  [1:0] v$3_32_out0;
wire  [1:0] v$6_998_out0;
wire  [1:0] v$6_999_out0;
wire  [1:0] v$8_112_out0;
wire  [1:0] v$8_113_out0;
wire  [1:0] v$9_1087_out0;
wire  [1:0] v$9_1088_out0;
wire  [1:0] v$AD1_5401_out0;
wire  [1:0] v$AD1_5402_out0;
wire  [1:0] v$AD2_4281_out0;
wire  [1:0] v$AD2_4282_out0;
wire  [1:0] v$AD3_4063_out0;
wire  [1:0] v$AD3_4064_out0;
wire  [1:0] v$C17_5068_out0;
wire  [1:0] v$C18_1516_out0;
wire  [1:0] v$C1_4009_out0;
wire  [1:0] v$C1_4010_out0;
wire  [1:0] v$C1_4681_out0;
wire  [1:0] v$C22_3079_out0;
wire  [1:0] v$C2_2749_out0;
wire  [1:0] v$C2_3117_out0;
wire  [1:0] v$C31_1111_out0;
wire  [1:0] v$C3_3893_out0;
wire  [1:0] v$C3_4484_out0;
wire  [1:0] v$C8_338_out0;
wire  [1:0] v$CONTROLREQUEST1_1141_out0;
wire  [1:0] v$CONTROLREQUEST2_4145_out0;
wire  [1:0] v$CONTROLREQUEST_2332_out0;
wire  [1:0] v$CONTROLREQUEST_2333_out0;
wire  [1:0] v$ControlRequest1_214_out0;
wire  [1:0] v$ControlRequest2_5031_out0;
wire  [1:0] v$D_2851_out0;
wire  [1:0] v$D_2852_out0;
wire  [1:0] v$D_5138_out0;
wire  [1:0] v$D_5139_out0;
wire  [1:0] v$D_539_out0;
wire  [1:0] v$D_540_out0;
wire  [1:0] v$INT_4565_out0;
wire  [1:0] v$MUX1_17_out0;
wire  [1:0] v$MUX1_18_out0;
wire  [1:0] v$MUX2_981_out0;
wire  [1:0] v$MUX2_982_out0;
wire  [1:0] v$M_1134_out0;
wire  [1:0] v$M_1135_out0;
wire  [1:0] v$M_4607_out0;
wire  [1:0] v$M_4608_out0;
wire  [1:0] v$NOTUSE2_4541_out0;
wire  [1:0] v$Q1_4523_out0;
wire  [1:0] v$Q1_4524_out0;
wire  [1:0] v$Q_3845_out0;
wire  [1:0] v$Q_3846_out0;
wire  [1:0] v$Q_5292_out0;
wire  [1:0] v$Q_5293_out0;
wire  [1:0] v$ROR_3251_out0;
wire  [1:0] v$ROR_3252_out0;
wire  [1:0] v$ROUNDING_3068_out0;
wire  [1:0] v$SEL2_817_out0;
wire  [1:0] v$SEL47_4498_out0;
wire  [1:0] v$SEL48_4857_out0;
wire  [1:0] v$SEL81_3767_out0;
wire  [1:0] v$SEL89_1033_out0;
wire  [1:0] v$SHIFTPREVIOUS_1586_out0;
wire  [1:0] v$SHIFTPREVIOUS_1587_out0;
wire  [1:0] v$SHIFT_1565_out0;
wire  [1:0] v$SHIFT_1566_out0;
wire  [1:0] v$SHIFT_2188_out0;
wire  [1:0] v$SHIFT_2189_out0;
wire  [1:0] v$SR_2469_out0;
wire  [1:0] v$SR_2470_out0;
wire  [1:0] v$SR_3148_out0;
wire  [1:0] v$SR_3149_out0;
wire  [1:0] v$SR_3994_out0;
wire  [1:0] v$SR_3995_out0;
wire  [1:0] v$SR_4135_out0;
wire  [1:0] v$SR_4136_out0;
wire  [1:0] v$SR_4826_out0;
wire  [1:0] v$SR_4827_out0;
wire  [1:0] v$SR_911_out0;
wire  [1:0] v$SR_912_out0;
wire  [1:0] v$X1_816_out0;
wire  [1:0] v$X8_2515_out0;
wire  [1:0] v$ZERO_3309_out0;
wire  [1:0] v$ZERO_3310_out0;
wire  [1:0] v$_1050_out0;
wire  [1:0] v$_1051_out0;
wire  [1:0] v$_1069_out0;
wire  [1:0] v$_1070_out0;
wire  [1:0] v$_1080_out1;
wire  [1:0] v$_1081_out1;
wire  [1:0] v$_1163_out0;
wire  [1:0] v$_1164_out0;
wire  [1:0] v$_1165_out0;
wire  [1:0] v$_1166_out0;
wire  [1:0] v$_116_out0;
wire  [1:0] v$_117_out0;
wire  [1:0] v$_118_out0;
wire  [1:0] v$_119_out0;
wire  [1:0] v$_120_out0;
wire  [1:0] v$_1212_out0;
wire  [1:0] v$_121_out0;
wire  [1:0] v$_122_out0;
wire  [1:0] v$_123_out0;
wire  [1:0] v$_124_out0;
wire  [1:0] v$_125_out0;
wire  [1:0] v$_126_out0;
wire  [1:0] v$_127_out0;
wire  [1:0] v$_128_out0;
wire  [1:0] v$_1430_out0;
wire  [1:0] v$_1431_out0;
wire  [1:0] v$_1432_out0;
wire  [1:0] v$_1433_out0;
wire  [1:0] v$_1562_out0;
wire  [1:0] v$_1607_out0;
wire  [1:0] v$_1608_out0;
wire  [1:0] v$_1609_out0;
wire  [1:0] v$_1610_out0;
wire  [1:0] v$_1660_out0;
wire  [1:0] v$_1661_out0;
wire  [1:0] v$_1720_out0;
wire  [1:0] v$_1721_out0;
wire  [1:0] v$_1723_out0;
wire  [1:0] v$_1746_out0;
wire  [1:0] v$_1747_out0;
wire  [1:0] v$_174_out0;
wire  [1:0] v$_175_out0;
wire  [1:0] v$_176_out0;
wire  [1:0] v$_1779_out0;
wire  [1:0] v$_177_out0;
wire  [1:0] v$_1797_out0;
wire  [1:0] v$_1809_out0;
wire  [1:0] v$_1878_out0;
wire  [1:0] v$_1888_out0;
wire  [1:0] v$_1889_out0;
wire  [1:0] v$_1890_out0;
wire  [1:0] v$_1891_out0;
wire  [1:0] v$_1912_out0;
wire  [1:0] v$_1913_out0;
wire  [1:0] v$_1914_out0;
wire  [1:0] v$_1915_out0;
wire  [1:0] v$_1916_out0;
wire  [1:0] v$_1917_out0;
wire  [1:0] v$_1918_out0;
wire  [1:0] v$_1919_out0;
wire  [1:0] v$_1920_out0;
wire  [1:0] v$_1921_out0;
wire  [1:0] v$_1922_out0;
wire  [1:0] v$_1965_out0;
wire  [1:0] v$_2097_out0;
wire  [1:0] v$_20_out0;
wire  [1:0] v$_2129_out0;
wire  [1:0] v$_21_out0;
wire  [1:0] v$_223_out1;
wire  [1:0] v$_224_out1;
wire  [1:0] v$_22_out0;
wire  [1:0] v$_2353_out0;
wire  [1:0] v$_2354_out0;
wire  [1:0] v$_2355_out0;
wire  [1:0] v$_2356_out0;
wire  [1:0] v$_236_out0;
wire  [1:0] v$_237_out0;
wire  [1:0] v$_238_out0;
wire  [1:0] v$_239_out0;
wire  [1:0] v$_2402_out0;
wire  [1:0] v$_2476_out0;
wire  [1:0] v$_2477_out0;
wire  [1:0] v$_2509_out0;
wire  [1:0] v$_2510_out0;
wire  [1:0] v$_2586_out1;
wire  [1:0] v$_2587_out1;
wire  [1:0] v$_2588_out1;
wire  [1:0] v$_2589_out1;
wire  [1:0] v$_2590_out1;
wire  [1:0] v$_2591_out1;
wire  [1:0] v$_2592_out1;
wire  [1:0] v$_2593_out1;
wire  [1:0] v$_2594_out1;
wire  [1:0] v$_2595_out1;
wire  [1:0] v$_2596_out1;
wire  [1:0] v$_2630_out0;
wire  [1:0] v$_2694_out0;
wire  [1:0] v$_2711_out0;
wire  [1:0] v$_2712_out0;
wire  [1:0] v$_2734_out0;
wire  [1:0] v$_2735_out0;
wire  [1:0] v$_2736_out0;
wire  [1:0] v$_2737_out0;
wire  [1:0] v$_2747_out1;
wire  [1:0] v$_2748_out1;
wire  [1:0] v$_2977_out0;
wire  [1:0] v$_2978_out0;
wire  [1:0] v$_2979_out0;
wire  [1:0] v$_2980_out0;
wire  [1:0] v$_3107_out0;
wire  [1:0] v$_3108_out0;
wire  [1:0] v$_3109_out0;
wire  [1:0] v$_3110_out0;
wire  [1:0] v$_3221_out0;
wire  [1:0] v$_3222_out0;
wire  [1:0] v$_3223_out0;
wire  [1:0] v$_3224_out0;
wire  [1:0] v$_3225_out0;
wire  [1:0] v$_3226_out0;
wire  [1:0] v$_3227_out0;
wire  [1:0] v$_3228_out0;
wire  [1:0] v$_3229_out0;
wire  [1:0] v$_3230_out0;
wire  [1:0] v$_3231_out0;
wire  [1:0] v$_3287_out0;
wire  [1:0] v$_3288_out0;
wire  [1:0] v$_3289_out0;
wire  [1:0] v$_3290_out0;
wire  [1:0] v$_3291_out0;
wire  [1:0] v$_3292_out0;
wire  [1:0] v$_3293_out0;
wire  [1:0] v$_3294_out0;
wire  [1:0] v$_3295_out0;
wire  [1:0] v$_3296_out0;
wire  [1:0] v$_3297_out0;
wire  [1:0] v$_3363_out0;
wire  [1:0] v$_3364_out0;
wire  [1:0] v$_3366_out0;
wire  [1:0] v$_3482_out0;
wire  [1:0] v$_3483_out0;
wire  [1:0] v$_3525_out1;
wire  [1:0] v$_3547_out0;
wire  [1:0] v$_3548_out0;
wire  [1:0] v$_3575_out0;
wire  [1:0] v$_3576_out0;
wire  [1:0] v$_3577_out0;
wire  [1:0] v$_3578_out0;
wire  [1:0] v$_3586_out0;
wire  [1:0] v$_3616_out0;
wire  [1:0] v$_3617_out0;
wire  [1:0] v$_361_out0;
wire  [1:0] v$_3624_out0;
wire  [1:0] v$_3625_out0;
wire  [1:0] v$_3626_out0;
wire  [1:0] v$_3627_out0;
wire  [1:0] v$_362_out0;
wire  [1:0] v$_3637_out0;
wire  [1:0] v$_3638_out0;
wire  [1:0] v$_3639_out0;
wire  [1:0] v$_363_out0;
wire  [1:0] v$_3640_out0;
wire  [1:0] v$_3710_out1;
wire  [1:0] v$_3814_out0;
wire  [1:0] v$_3815_out0;
wire  [1:0] v$_3816_out0;
wire  [1:0] v$_3817_out0;
wire  [1:0] v$_3877_out0;
wire  [1:0] v$_3878_out0;
wire  [1:0] v$_404_out0;
wire  [1:0] v$_4073_out0;
wire  [1:0] v$_4126_out0;
wire  [1:0] v$_4127_out0;
wire  [1:0] v$_4128_out0;
wire  [1:0] v$_4129_out0;
wire  [1:0] v$_4258_out0;
wire  [1:0] v$_4259_out0;
wire  [1:0] v$_4270_out0;
wire  [1:0] v$_4271_out0;
wire  [1:0] v$_4408_out0;
wire  [1:0] v$_4409_out0;
wire  [1:0] v$_4438_out0;
wire  [1:0] v$_4491_out0;
wire  [1:0] v$_4662_out0;
wire  [1:0] v$_4663_out0;
wire  [1:0] v$_4664_out0;
wire  [1:0] v$_4665_out0;
wire  [1:0] v$_4666_out0;
wire  [1:0] v$_4667_out0;
wire  [1:0] v$_4668_out0;
wire  [1:0] v$_4669_out0;
wire  [1:0] v$_4670_out0;
wire  [1:0] v$_4671_out0;
wire  [1:0] v$_4672_out0;
wire  [1:0] v$_4769_out0;
wire  [1:0] v$_4788_out0;
wire  [1:0] v$_4789_out0;
wire  [1:0] v$_4790_out0;
wire  [1:0] v$_483_out0;
wire  [1:0] v$_484_out0;
wire  [1:0] v$_4858_out0;
wire  [1:0] v$_485_out0;
wire  [1:0] v$_4862_out0;
wire  [1:0] v$_4878_out0;
wire  [1:0] v$_4879_out0;
wire  [1:0] v$_4880_out0;
wire  [1:0] v$_4881_out0;
wire  [1:0] v$_4938_out1;
wire  [1:0] v$_4968_out0;
wire  [1:0] v$_4969_out0;
wire  [1:0] v$_498_out0;
wire  [1:0] v$_5136_out0;
wire  [1:0] v$_5137_out0;
wire  [1:0] v$_5259_out0;
wire  [1:0] v$_5414_out0;
wire  [1:0] v$_5415_out0;
wire  [1:0] v$_717_out0;
wire  [1:0] v$_773_out1;
wire  [1:0] v$_774_out1;
wire  [1:0] v$_839_out0;
wire  [1:0] v$_840_out0;
wire  [1:0] v$_841_out0;
wire  [1:0] v$_842_out0;
wire  [1:0] v$_943_out0;
wire  [1:0] v$_944_out0;
wire  [1:0] v$_945_out0;
wire  [1:0] v$_946_out0;
wire  [20:0] v$00_1369_out0;
wire  [20:0] v$1_4825_out0;
wire  [20:0] v$B10_317_out0;
wire  [20:0] v$B10_4097_out0;
wire  [20:0] v$MUX11_990_out0;
wire  [20:0] v$MUX12_4386_out0;
wire  [20:0] v$MUX13_300_out0;
wire  [20:0] v$MUX18_2756_out0;
wire  [20:0] v$MUX1_533_out0;
wire  [20:0] v$MUX20_5281_out0;
wire  [20:0] v$MUX21_762_out0;
wire  [20:0] v$MUX23_3043_out0;
wire  [20:0] v$MUX24_3282_out0;
wire  [20:0] v$MUX25_1038_out0;
wire  [20:0] v$MUX27_2678_out0;
wire  [20:0] v$MUX28_5060_out0;
wire  [20:0] v$MUX2_3635_out0;
wire  [20:0] v$MUX3_5301_out0;
wire  [20:0] v$MUX4_3788_out0;
wire  [20:0] v$MUX5_3531_out0;
wire  [20:0] v$MUX6_5312_out0;
wire  [20:0] v$MUX7_1475_out0;
wire  [20:0] v$MUX8_1156_out0;
wire  [20:0] v$MUX9_2441_out0;
wire  [20:0] v$N2_2836_out0;
wire  [20:0] v$N2_680_out0;
wire  [20:0] v$N2_820_out0;
wire  [20:0] v$N3_3326_out0;
wire  [20:0] v$N3_3728_out0;
wire  [20:0] v$N3_4935_out0;
wire  [20:0] v$OUTPUT_5043_out0;
wire  [20:0] v$_0_out0;
wire  [20:0] v$_1099_out0;
wire  [20:0] v$_10_out0;
wire  [20:0] v$_1241_out0;
wire  [20:0] v$_1264_out0;
wire  [20:0] v$_1906_out0;
wire  [20:0] v$_2006_out0;
wire  [20:0] v$_2131_out0;
wire  [20:0] v$_2422_out0;
wire  [20:0] v$_2865_out0;
wire  [20:0] v$_3128_out0;
wire  [20:0] v$_3261_out0;
wire  [20:0] v$_3335_out1;
wire  [20:0] v$_33_out0;
wire  [20:0] v$_416_out0;
wire  [20:0] v$_4209_out0;
wire  [20:0] v$_4415_out0;
wire  [20:0] v$_4446_out0;
wire  [20:0] v$_4647_out0;
wire  [20:0] v$_4773_out0;
wire  [20:0] v$_5032_out0;
wire  [20:0] v$_5096_out1;
wire  [20:0] v$_5220_out0;
wire  [20:0] v$_5245_out0;
wire  [20:0] v$_5248_out0;
wire  [20:0] v$_5389_out0;
wire  [20:0] v$_5424_out0;
wire  [20:0] v$_588_out0;
wire  [20:0] v$_635_out0;
wire  [20:0] v$_708_out0;
wire  [20:0] v$_728_out0;
wire  [20:0] v$_980_out0;
wire  [21:0] v$11_2653_out0;
wire  [21:0] v$FRAC22_4051_out0;
wire  [21:0] v$FRAC_1303_out0;
wire  [21:0] v$IN1_3927_out0;
wire  [21:0] v$INPUT_2972_out0;
wire  [21:0] v$IN_1444_out0;
wire  [21:0] v$MUX10_1398_out0;
wire  [21:0] v$MUX11_3385_out0;
wire  [21:0] v$MUX12_4718_out0;
wire  [21:0] v$MUX2_5410_out0;
wire  [21:0] v$MUX2_974_out0;
wire  [21:0] v$MUX3_1699_out0;
wire  [21:0] v$MUX3_4210_out0;
wire  [21:0] v$MUX4_3839_out0;
wire  [21:0] v$MUX4_48_out0;
wire  [21:0] v$MUX5_156_out0;
wire  [21:0] v$MUX6_1531_out0;
wire  [21:0] v$MUX7_4758_out0;
wire  [21:0] v$MUX8_349_out0;
wire  [21:0] v$MUX9_3900_out0;
wire  [21:0] v$NEWFRAC0001_4382_out0;
wire  [21:0] v$NEWFRAC1011_2046_out0;
wire  [21:0] v$NEWFRAC_249_out0;
wire  [21:0] v$OUT1_1685_out0;
wire  [21:0] v$OUTPUT_1902_out0;
wire  [21:0] v$OUT_3656_out0;
wire  [21:0] v$_1417_out0;
wire  [21:0] v$_157_out0;
wire  [21:0] v$_1735_out0;
wire  [21:0] v$_2181_out0;
wire  [21:0] v$_2375_out0;
wire  [21:0] v$_2456_out0;
wire  [21:0] v$_2772_out0;
wire  [21:0] v$_2838_out0;
wire  [21:0] v$_2849_out0;
wire  [21:0] v$_3708_out0;
wire  [21:0] v$_3724_out0;
wire  [21:0] v$_3926_out0;
wire  [21:0] v$_4616_out0;
wire  [21:0] v$_5250_out0;
wire  [21:0] v$_58_out0;
wire  [21:0] v$_716_out0;
wire  [22:0] v$_350_out0;
wire  [23:0] v$_942_out0;
wire  [27:0] v$_3365_out0;
wire  [27:0] v$_5115_out0;
wire  [27:0] v$_5116_out0;
wire  [28:0] v$CONTROLPROTOCAL1_4086_out0;
wire  [28:0] v$CONTROLPROTOCAL2_1243_out0;
wire  [28:0] v$MUX1_2742_out0;
wire  [28:0] v$WEN$DATA1_3913_out0;
wire  [28:0] v$WEN$DATA2_3530_out0;
wire  [28:0] v$WENDATA1_1446_out0;
wire  [28:0] v$WENDATA2_2308_out0;
wire  [28:0] v$WENDATA_162_out0;
wire  [28:0] v$WENDATA_163_out0;
wire  [28:0] v$_2654_out0;
wire  [28:0] v$_2655_out0;
wire  [2:0] v$1_4387_out0;
wire  [2:0] v$1_4388_out0;
wire  [2:0] v$C18_1515_out0;
wire  [2:0] v$C3_3005_out0;
wire  [2:0] v$C3_4571_out0;
wire  [2:0] v$C3_4882_out0;
wire  [2:0] v$C4_2077_out0;
wire  [2:0] v$C4_627_out0;
wire  [2:0] v$C6_3912_out0;
wire  [2:0] v$NA_3557_out0;
wire  [2:0] v$NA_3558_out0;
wire  [2:0] v$OP_534_out0;
wire  [2:0] v$OP_535_out0;
wire  [2:0] v$OP_966_out0;
wire  [2:0] v$OP_967_out0;
wire  [2:0] v$SEL68_3726_out0;
wire  [2:0] v$X2_531_out0;
wire  [2:0] v$X6_673_out0;
wire  [2:0] v$_1178_out0;
wire  [2:0] v$_1179_out0;
wire  [2:0] v$_1180_out0;
wire  [2:0] v$_1386_out0;
wire  [2:0] v$_1419_out0;
wire  [2:0] v$_1593_out0;
wire  [2:0] v$_2111_out1;
wire  [2:0] v$_2112_out1;
wire  [2:0] v$_2113_out1;
wire  [2:0] v$_2114_out1;
wire  [2:0] v$_2115_out1;
wire  [2:0] v$_2116_out1;
wire  [2:0] v$_2117_out1;
wire  [2:0] v$_2118_out1;
wire  [2:0] v$_2119_out1;
wire  [2:0] v$_2120_out1;
wire  [2:0] v$_2121_out1;
wire  [2:0] v$_2428_out0;
wire  [2:0] v$_2926_out0;
wire  [2:0] v$_2949_out1;
wire  [2:0] v$_2950_out1;
wire  [2:0] v$_3121_out0;
wire  [2:0] v$_3618_out1;
wire  [2:0] v$_3677_out0;
wire  [2:0] v$_4804_out1;
wire  [2:0] v$_4805_out1;
wire  [2:0] v$_5062_out0;
wire  [2:0] v$_5063_out0;
wire  [2:0] v$_5317_out1;
wire  [2:0] v$_5318_out1;
wire  [2:0] v$_532_out0;
wire  [2:0] v$_5433_out0;
wire  [2:0] v$_5434_out0;
wire  [2:0] v$_5435_out0;
wire  [2:0] v$_5436_out0;
wire  [2:0] v$_5437_out0;
wire  [2:0] v$_5438_out0;
wire  [2:0] v$_5439_out0;
wire  [2:0] v$_5440_out0;
wire  [2:0] v$_5441_out0;
wire  [2:0] v$_5442_out0;
wire  [2:0] v$_5443_out0;
wire  [2:0] v$_776_out0;
wire  [2:0] v$_972_out0;
wire  [3:0] v$4_2287_out0;
wire  [3:0] v$4_2288_out0;
wire  [3:0] v$5_609_out0;
wire  [3:0] v$5_610_out0;
wire  [3:0] v$9_3069_out0;
wire  [3:0] v$9_3070_out0;
wire  [3:0] v$B_1966_out0;
wire  [3:0] v$B_1967_out0;
wire  [3:0] v$B_3493_out0;
wire  [3:0] v$B_3494_out0;
wire  [3:0] v$B_578_out0;
wire  [3:0] v$B_579_out0;
wire  [3:0] v$B_985_out0;
wire  [3:0] v$B_986_out0;
wire  [3:0] v$C10_1253_out0;
wire  [3:0] v$C10_1968_out0;
wire  [3:0] v$C10_1969_out0;
wire  [3:0] v$C11_3342_out0;
wire  [3:0] v$C11_3343_out0;
wire  [3:0] v$C11_3383_out0;
wire  [3:0] v$C12_2310_out0;
wire  [3:0] v$C12_2311_out0;
wire  [3:0] v$C13_1292_out0;
wire  [3:0] v$C13_1293_out0;
wire  [3:0] v$C14_2740_out0;
wire  [3:0] v$C14_2741_out0;
wire  [3:0] v$C1_2298_out0;
wire  [3:0] v$C1_2299_out0;
wire  [3:0] v$C1_3658_out0;
wire  [3:0] v$C1_3659_out0;
wire  [3:0] v$C26_1186_out0;
wire  [3:0] v$C2_4459_out0;
wire  [3:0] v$C2_4460_out0;
wire  [3:0] v$C3_5357_out0;
wire  [3:0] v$C3_5358_out0;
wire  [3:0] v$C4_1031_out0;
wire  [3:0] v$C4_1032_out0;
wire  [3:0] v$C4_2007_out0;
wire  [3:0] v$C5_1899_out0;
wire  [3:0] v$C5_4214_out0;
wire  [3:0] v$C5_4464_out0;
wire  [3:0] v$C5_4465_out0;
wire  [3:0] v$C6_4823_out0;
wire  [3:0] v$C6_4824_out0;
wire  [3:0] v$C7_1908_out0;
wire  [3:0] v$C7_1909_out0;
wire  [3:0] v$C8_2634_out0;
wire  [3:0] v$C8_2635_out0;
wire  [3:0] v$C9_2796_out0;
wire  [3:0] v$C9_2797_out0;
wire  [3:0] v$MUX10_589_out0;
wire  [3:0] v$MUX10_590_out0;
wire  [3:0] v$MUX11_1881_out0;
wire  [3:0] v$MUX11_1882_out0;
wire  [3:0] v$MUX12_3905_out0;
wire  [3:0] v$MUX12_3906_out0;
wire  [3:0] v$MUX13_849_out0;
wire  [3:0] v$MUX13_850_out0;
wire  [3:0] v$MUX1_2932_out0;
wire  [3:0] v$MUX1_2933_out0;
wire  [3:0] v$MUX2_1039_out0;
wire  [3:0] v$MUX2_1040_out0;
wire  [3:0] v$MUX3_2997_out0;
wire  [3:0] v$MUX3_2998_out0;
wire  [3:0] v$MUX4_725_out0;
wire  [3:0] v$MUX4_726_out0;
wire  [3:0] v$MUX5_1751_out0;
wire  [3:0] v$MUX5_1752_out0;
wire  [3:0] v$MUX6_3118_out0;
wire  [3:0] v$MUX6_3119_out0;
wire  [3:0] v$MUX7_525_out0;
wire  [3:0] v$MUX7_526_out0;
wire  [3:0] v$MUX8_2408_out0;
wire  [3:0] v$MUX8_2409_out0;
wire  [3:0] v$MUX9_3445_out0;
wire  [3:0] v$MUX9_3446_out0;
wire  [3:0] v$NOTUSE4_5218_out0;
wire  [3:0] v$NOTUSED_4762_out0;
wire  [3:0] v$NOTUSED_4763_out0;
wire  [3:0] v$NOTUSE_2579_out0;
wire  [3:0] v$N_2709_out0;
wire  [3:0] v$N_2710_out0;
wire  [3:0] v$N_5197_out0;
wire  [3:0] v$N_5198_out0;
wire  [3:0] v$O_2429_out0;
wire  [3:0] v$O_2430_out0;
wire  [3:0] v$SEL1_565_out0;
wire  [3:0] v$SEL1_566_out0;
wire  [3:0] v$SEL7_3629_out0;
wire  [3:0] v$SHIFTNUMBER_336_out0;
wire  [3:0] v$SHIFTNUMBER_337_out0;
wire  [3:0] v$SHIFTNUMBER_5177_out0;
wire  [3:0] v$X11_3193_out0;
wire  [3:0] v$X3_1541_out0;
wire  [3:0] v$ZERO_3207_out0;
wire  [3:0] v$ZERO_3208_out0;
wire  [3:0] v$_1001_out0;
wire  [3:0] v$_1002_out0;
wire  [3:0] v$_1003_out0;
wire  [3:0] v$_1297_out1;
wire  [3:0] v$_1298_out1;
wire  [3:0] v$_1320_out0;
wire  [3:0] v$_1420_out0;
wire  [3:0] v$_1421_out0;
wire  [3:0] v$_1422_out0;
wire  [3:0] v$_1423_out0;
wire  [3:0] v$_1527_out0;
wire  [3:0] v$_1528_out0;
wire  [3:0] v$_1603_out0;
wire  [3:0] v$_1604_out0;
wire  [3:0] v$_1605_out0;
wire  [3:0] v$_1606_out0;
wire  [3:0] v$_1670_out0;
wire  [3:0] v$_1671_out0;
wire  [3:0] v$_1672_out0;
wire  [3:0] v$_1673_out0;
wire  [3:0] v$_1940_out0;
wire  [3:0] v$_1941_out0;
wire  [3:0] v$_1942_out0;
wire  [3:0] v$_1943_out0;
wire  [3:0] v$_1944_out0;
wire  [3:0] v$_1945_out0;
wire  [3:0] v$_1946_out0;
wire  [3:0] v$_1947_out0;
wire  [3:0] v$_1948_out0;
wire  [3:0] v$_1949_out0;
wire  [3:0] v$_1950_out0;
wire  [3:0] v$_2017_out0;
wire  [3:0] v$_2018_out0;
wire  [3:0] v$_2019_out0;
wire  [3:0] v$_2020_out0;
wire  [3:0] v$_2073_out0;
wire  [3:0] v$_2074_out0;
wire  [3:0] v$_2075_out0;
wire  [3:0] v$_2076_out0;
wire  [3:0] v$_2148_out1;
wire  [3:0] v$_2149_out1;
wire  [3:0] v$_2150_out1;
wire  [3:0] v$_2151_out1;
wire  [3:0] v$_2152_out1;
wire  [3:0] v$_2153_out1;
wire  [3:0] v$_2154_out1;
wire  [3:0] v$_2155_out1;
wire  [3:0] v$_2156_out1;
wire  [3:0] v$_2157_out1;
wire  [3:0] v$_2158_out1;
wire  [3:0] v$_2192_out0;
wire  [3:0] v$_2328_out0;
wire  [3:0] v$_2329_out0;
wire  [3:0] v$_2342_out0;
wire  [3:0] v$_2343_out0;
wire  [3:0] v$_2344_out0;
wire  [3:0] v$_2345_out0;
wire  [3:0] v$_2346_out0;
wire  [3:0] v$_2347_out0;
wire  [3:0] v$_2348_out0;
wire  [3:0] v$_2349_out0;
wire  [3:0] v$_2350_out0;
wire  [3:0] v$_2351_out0;
wire  [3:0] v$_2352_out0;
wire  [3:0] v$_2620_out0;
wire  [3:0] v$_2621_out0;
wire  [3:0] v$_2623_out1;
wire  [3:0] v$_2624_out1;
wire  [3:0] v$_2658_out0;
wire  [3:0] v$_2659_out0;
wire  [3:0] v$_2660_out0;
wire  [3:0] v$_2661_out0;
wire  [3:0] v$_2705_out0;
wire  [3:0] v$_272_out0;
wire  [3:0] v$_2787_out0;
wire  [3:0] v$_2788_out0;
wire  [3:0] v$_3120_out0;
wire  [3:0] v$_3122_out0;
wire  [3:0] v$_316_out0;
wire  [3:0] v$_3346_out1;
wire  [3:0] v$_3347_out1;
wire  [3:0] v$_3422_out1;
wire  [3:0] v$_3423_out1;
wire  [3:0] v$_3591_out0;
wire  [3:0] v$_3592_out0;
wire  [3:0] v$_3599_out0;
wire  [3:0] v$_3600_out0;
wire  [3:0] v$_3621_out0;
wire  [3:0] v$_3622_out0;
wire  [3:0] v$_3623_out0;
wire  [3:0] v$_365_out0;
wire  [3:0] v$_3725_out0;
wire  [3:0] v$_3740_out1;
wire  [3:0] v$_376_out0;
wire  [3:0] v$_399_out0;
wire  [3:0] v$_400_out0;
wire  [3:0] v$_4157_out0;
wire  [3:0] v$_4158_out0;
wire  [3:0] v$_4159_out0;
wire  [3:0] v$_4160_out0;
wire  [3:0] v$_4393_out0;
wire  [3:0] v$_4475_out0;
wire  [3:0] v$_4504_out1;
wire  [3:0] v$_4505_out1;
wire  [3:0] v$_4717_out0;
wire  [3:0] v$_4753_out0;
wire  [3:0] v$_4754_out0;
wire  [3:0] v$_4755_out0;
wire  [3:0] v$_4756_out0;
wire  [3:0] v$_4766_out1;
wire  [3:0] v$_4870_out0;
wire  [3:0] v$_5276_out0;
wire  [3:0] v$_5277_out0;
wire  [4:0] v$4_2262_out0;
wire  [4:0] v$4_2263_out0;
wire  [4:0] v$A1_1910_out0;
wire  [4:0] v$A1_5395_out0;
wire  [4:0] v$A2_528_out0;
wire  [4:0] v$BIGGEREXPO_1814_out0;
wire  [4:0] v$C10_2986_out0;
wire  [4:0] v$C10_3628_out0;
wire  [4:0] v$C11_3973_out0;
wire  [4:0] v$C12_1322_out0;
wire  [4:0] v$C13_5266_out0;
wire  [4:0] v$C14_576_out0;
wire  [4:0] v$C15_2147_out0;
wire  [4:0] v$C16_205_out0;
wire  [4:0] v$C16_206_out0;
wire  [4:0] v$C16_427_out0;
wire  [4:0] v$C17_1139_out0;
wire  [4:0] v$C17_5302_out0;
wire  [4:0] v$C18_3898_out0;
wire  [4:0] v$C19_5406_out0;
wire  [4:0] v$C1_2206_out0;
wire  [4:0] v$C1_2374_out0;
wire  [4:0] v$C1_2666_out0;
wire  [4:0] v$C1_4327_out0;
wire  [4:0] v$C20_1438_out0;
wire  [4:0] v$C20_4877_out0;
wire  [4:0] v$C21_5199_out0;
wire  [4:0] v$C22_372_out0;
wire  [4:0] v$C27_3680_out0;
wire  [4:0] v$C28_1010_out0;
wire  [4:0] v$C28_1203_out0;
wire  [4:0] v$C2_2234_out0;
wire  [4:0] v$C2_3555_out0;
wire  [4:0] v$C30_4304_out0;
wire  [4:0] v$C30_536_out0;
wire  [4:0] v$C31_3551_out0;
wire  [4:0] v$C3_1385_out0;
wire  [4:0] v$C4_3256_out0;
wire  [4:0] v$C4_777_out0;
wire  [4:0] v$C5_4307_out0;
wire  [4:0] v$C6_2426_out0;
wire  [4:0] v$C6_3198_out0;
wire  [4:0] v$C6_3481_out0;
wire  [4:0] v$C6_34_out0;
wire  [4:0] v$C7_2066_out0;
wire  [4:0] v$C8_13_out0;
wire  [4:0] v$C8_3052_out0;
wire  [4:0] v$C9_1415_out0;
wire  [4:0] v$C9_3886_out0;
wire  [4:0] v$DIFFERENCE_133_out0;
wire  [4:0] v$DIFFERENCE_5352_out0;
wire  [4:0] v$EXPA_1502_out0;
wire  [4:0] v$EXPA_4353_out0;
wire  [4:0] v$EXPB_3248_out0;
wire  [4:0] v$EXPB_3876_out0;
wire  [4:0] v$EXPO0IFNEG_1045_out0;
wire  [4:0] v$EXPOA_1226_out0;
wire  [4:0] v$EXPOA_1813_out0;
wire  [4:0] v$EXPOA_2078_out0;
wire  [4:0] v$EXPOB_1579_out0;
wire  [4:0] v$EXPOB_3402_out0;
wire  [4:0] v$EXPOB_5159_out0;
wire  [4:0] v$EXPODIFF_3582_out0;
wire  [4:0] v$EXPODIFF_4412_out0;
wire  [4:0] v$EXPONENTA_1574_out0;
wire  [4:0] v$EXPONENTB_2080_out0;
wire  [4:0] v$EXPONENTDIFFERENCE13_2330_out0;
wire  [4:0] v$EXPONENT_245_out0;
wire  [4:0] v$EXPONENT_2696_out0;
wire  [4:0] v$EXPONENT_4661_out0;
wire  [4:0] v$EXPONENT_5291_out0;
wire  [4:0] v$EXPONENT_95_out0;
wire  [4:0] v$K_135_out0;
wire  [4:0] v$K_136_out0;
wire  [4:0] v$MUX11_5024_out0;
wire  [4:0] v$MUX12_4936_out0;
wire  [4:0] v$MUX13_1767_out0;
wire  [4:0] v$MUX14_142_out0;
wire  [4:0] v$MUX14_3139_out0;
wire  [4:0] v$MUX15_1450_out0;
wire  [4:0] v$MUX15_5222_out0;
wire  [4:0] v$MUX15_5223_out0;
wire  [4:0] v$MUX16_4015_out0;
wire  [4:0] v$MUX16_907_out0;
wire  [4:0] v$MUX16_908_out0;
wire  [4:0] v$MUX17_3354_out0;
wire  [4:0] v$MUX18_5418_out0;
wire  [4:0] v$MUX19_2194_out0;
wire  [4:0] v$MUX1_3829_out0;
wire  [4:0] v$MUX1_493_out0;
wire  [4:0] v$MUX20_4105_out0;
wire  [4:0] v$MUX21_3934_out0;
wire  [4:0] v$MUX22_3031_out0;
wire  [4:0] v$MUX22_5423_out0;
wire  [4:0] v$MUX23_5205_out0;
wire  [4:0] v$MUX25_5182_out0;
wire  [4:0] v$MUX28_810_out0;
wire  [4:0] v$MUX2_37_out0;
wire  [4:0] v$MUX2_5303_out0;
wire  [4:0] v$MUX31_1588_out0;
wire  [4:0] v$MUX3_2558_out0;
wire  [4:0] v$MUX3_4060_out0;
wire  [4:0] v$MUX3_527_out0;
wire  [4:0] v$MUX4_1182_out0;
wire  [4:0] v$MUX4_4779_out0;
wire  [4:0] v$MUX4_5413_out0;
wire  [4:0] v$MUX5_1030_out0;
wire  [4:0] v$MUX5_3998_out0;
wire  [4:0] v$MUX6_3257_out0;
wire  [4:0] v$MUX7_685_out0;
wire  [4:0] v$MUX8_4023_out0;
wire  [4:0] v$NEWEXPO0001_1724_out0;
wire  [4:0] v$NEWEXPO1011_4381_out0;
wire  [4:0] v$NEWEXPONENT_1710_out0;
wire  [4:0] v$NEWEXPONENT_1711_out0;
wire  [4:0] v$NEWEXPO_4385_out0;
wire  [4:0] v$NEWEXPO_4492_out0;
wire  [4:0] v$NEWEXPO_5072_out0;
wire  [4:0] v$SEL1_1118_out0;
wire  [4:0] v$SEL1_3647_out0;
wire  [4:0] v$SEL2_3828_out0;
wire  [4:0] v$SEL2_814_out0;
wire  [4:0] v$SEL41_975_out0;
wire  [4:0] v$SEL4_1457_out0;
wire  [4:0] v$SEL6_3327_out0;
wire  [4:0] v$SHIFTNUMBER1_611_out0;
wire  [4:0] v$SHIFTNUMBER5_3520_out0;
wire  [4:0] v$SHIFTNUMBER_3013_out0;
wire  [4:0] v$SHIFTNUMBER_3952_out0;
wire  [4:0] v$SHIFTNUMBER_5176_out0;
wire  [4:0] v$SHIFTNUMBER_672_out0;
wire  [4:0] v$SHIFTNUM_5219_out0;
wire  [4:0] v$X2_3685_out0;
wire  [4:0] v$X5_134_out0;
wire  [4:0] v$XOR1_16_out0;
wire  [4:0] v$XOR2_5112_out0;
wire  [4:0] v$_1046_out0;
wire  [4:0] v$_1871_out0;
wire  [4:0] v$_2089_out1;
wire  [4:0] v$_242_out1;
wire  [4:0] v$_243_out1;
wire  [4:0] v$_2462_out0;
wire  [4:0] v$_2463_out0;
wire  [4:0] v$_2464_out0;
wire  [4:0] v$_2465_out0;
wire  [4:0] v$_3035_out0;
wire  [4:0] v$_3066_out0;
wire  [4:0] v$_3372_out0;
wire  [4:0] v$_3605_out0;
wire  [4:0] v$_3606_out0;
wire  [4:0] v$_3607_out0;
wire  [4:0] v$_4322_out0;
wire  [4:0] v$_4323_out0;
wire  [4:0] v$_4324_out0;
wire  [4:0] v$_4325_out0;
wire  [4:0] v$_4420_out1;
wire  [4:0] v$_4421_out1;
wire  [4:0] v$_4422_out1;
wire  [4:0] v$_4423_out1;
wire  [4:0] v$_4424_out1;
wire  [4:0] v$_4425_out1;
wire  [4:0] v$_4426_out1;
wire  [4:0] v$_4427_out1;
wire  [4:0] v$_4428_out1;
wire  [4:0] v$_4429_out1;
wire  [4:0] v$_4430_out1;
wire  [4:0] v$_4449_out0;
wire  [4:0] v$_4450_out0;
wire  [4:0] v$_4451_out0;
wire  [4:0] v$_4542_out0;
wire  [4:0] v$_4653_out0;
wire  [4:0] v$_4691_out0;
wire  [4:0] v$_5027_out1;
wire  [4:0] v$_5028_out1;
wire  [4:0] v$_863_out0;
wire  [4:0] v$comparator_4432_out0;
wire  [5:0] v$A1_2126_out0;
wire  [5:0] v$A1_2427_out0;
wire  [5:0] v$C15_3897_out0;
wire  [5:0] v$C1_3138_out0;
wire  [5:0] v$C2_3735_out0;
wire  [5:0] v$C5_2191_out0;
wire  [5:0] v$C5_4278_out0;
wire  [5:0] v$C6_3524_out0;
wire  [5:0] v$C6_5119_out0;
wire  [5:0] v$C7_228_out0;
wire  [5:0] v$MUX1_2143_out0;
wire  [5:0] v$SEL4_676_out0;
wire  [5:0] v$SEL51_4277_out0;
wire  [5:0] v$X15_2619_out0;
wire  [5:0] v$X4_3285_out0;
wire  [5:0] v$XOR1_3486_out0;
wire  [5:0] v$_1209_out0;
wire  [5:0] v$_1210_out0;
wire  [5:0] v$_1211_out0;
wire  [5:0] v$_1688_out0;
wire  [5:0] v$_1812_out0;
wire  [5:0] v$_2024_out0;
wire  [5:0] v$_2717_out1;
wire  [5:0] v$_2718_out1;
wire  [5:0] v$_3087_out0;
wire  [5:0] v$_3583_out0;
wire  [5:0] v$_4056_out0;
wire  [5:0] v$_4057_out0;
wire  [5:0] v$_4058_out0;
wire  [5:0] v$_4059_out0;
wire  [5:0] v$_4372_out1;
wire  [5:0] v$_4633_out1;
wire  [5:0] v$_4634_out1;
wire  [5:0] v$_4749_out0;
wire  [5:0] v$_482_out0;
wire  [5:0] v$_4832_out1;
wire  [5:0] v$_4833_out1;
wire  [5:0] v$_4834_out1;
wire  [5:0] v$_4835_out1;
wire  [5:0] v$_4836_out1;
wire  [5:0] v$_4837_out1;
wire  [5:0] v$_4838_out1;
wire  [5:0] v$_4839_out1;
wire  [5:0] v$_4840_out1;
wire  [5:0] v$_4841_out1;
wire  [5:0] v$_4842_out1;
wire  [5:0] v$_5167_out0;
wire  [5:0] v$_5278_out0;
wire  [5:0] v$_687_out0;
wire  [5:0] v$_688_out0;
wire  [5:0] v$_689_out0;
wire  [5:0] v$_690_out0;
wire  [5:0] v$_836_out0;
wire  [6:0] v$$EXPONENT_225_out0;
wire  [6:0] v$A1_2039_out0;
wire  [6:0] v$A2_4445_out0;
wire  [6:0] v$ABSOLUTE_486_out0;
wire  [6:0] v$C10_2703_out0;
wire  [6:0] v$C13_1573_out0;
wire  [6:0] v$C13_274_out0;
wire  [6:0] v$C15_4273_out0;
wire  [6:0] v$C2_4547_out0;
wire  [6:0] v$C7_5237_out0;
wire  [6:0] v$C7_825_out0;
wire  [6:0] v$C8_4082_out0;
wire  [6:0] v$C9_4326_out0;
wire  [6:0] v$DIFFERENCE7_132_out0;
wire  [6:0] v$EXPONENT_5089_out0;
wire  [6:0] v$EXPONENT_5290_out0;
wire  [6:0] v$EXPONENT_5297_out0;
wire  [6:0] v$EXPO_2336_out0;
wire  [6:0] v$EXPO_44_out0;
wire  [6:0] v$MUX14_141_out0;
wire  [6:0] v$NA_1621_out0;
wire  [6:0] v$NA_1622_out0;
wire  [6:0] v$SHIFT_3099_out0;
wire  [6:0] v$X22_2650_out0;
wire  [6:0] v$X7_4476_out0;
wire  [6:0] v$XOR1_1741_out0;
wire  [6:0] v$_1127_out0;
wire  [6:0] v$_159_out0;
wire  [6:0] v$_160_out0;
wire  [6:0] v$_161_out0;
wire  [6:0] v$_1903_out0;
wire  [6:0] v$_2639_out0;
wire  [6:0] v$_2649_out0;
wire  [6:0] v$_2760_out1;
wire  [6:0] v$_2761_out1;
wire  [6:0] v$_3090_out1;
wire  [6:0] v$_3556_out0;
wire  [6:0] v$_3745_out1;
wire  [6:0] v$_3746_out1;
wire  [6:0] v$_3747_out1;
wire  [6:0] v$_3748_out1;
wire  [6:0] v$_3749_out1;
wire  [6:0] v$_3750_out1;
wire  [6:0] v$_3751_out1;
wire  [6:0] v$_3752_out1;
wire  [6:0] v$_3753_out1;
wire  [6:0] v$_3754_out1;
wire  [6:0] v$_3755_out1;
wire  [6:0] v$_3832_out0;
wire  [6:0] v$_3833_out0;
wire  [6:0] v$_4095_out0;
wire  [6:0] v$_4250_out1;
wire  [6:0] v$_4251_out1;
wire  [6:0] v$_4863_out0;
wire  [6:0] v$_5429_out0;
wire  [6:0] v$_862_out0;
wire  [7:0] v$15TO8_5054_out0;
wire  [7:0] v$15TO8_5055_out0;
wire  [7:0] v$7TO0_3572_out0;
wire  [7:0] v$7TO0_3573_out0;
wire  [7:0] v$A1_2125_out0;
wire  [7:0] v$A_4699_out0;
wire  [7:0] v$B_2057_out0;
wire  [7:0] v$C15_3896_out0;
wire  [7:0] v$C1_2376_out0;
wire  [7:0] v$C1_2377_out0;
wire  [7:0] v$C24_2887_out0;
wire  [7:0] v$C4_1537_out0;
wire  [7:0] v$C5_4673_out0;
wire  [7:0] v$C8_4137_out0;
wire  [7:0] v$C8_598_out0;
wire  [7:0] v$C9_758_out0;
wire  [7:0] v$C_2732_out0;
wire  [7:0] v$INPUT_3072_out0;
wire  [7:0] v$NOTUSE2_3657_out0;
wire  [7:0] v$NOTUSE8_4490_out0;
wire  [7:0] v$OUTPUTSHIFT_5150_out0;
wire  [7:0] v$OUTPUT_1820_out0;
wire  [7:0] v$S1_2964_out0;
wire  [7:0] v$S2_2248_out0;
wire  [7:0] v$SEL49_3044_out0;
wire  [7:0] v$SEL51_2334_out0;
wire  [7:0] v$SEL52_902_out0;
wire  [7:0] v$X4_4257_out0;
wire  [7:0] v$X6_230_out0;
wire  [7:0] v$XOR1_3485_out0;
wire  [7:0] v$ZERO_295_out0;
wire  [7:0] v$ZERO_296_out0;
wire  [7:0] v$_1278_out1;
wire  [7:0] v$_1323_out0;
wire  [7:0] v$_1387_out0;
wire  [7:0] v$_14_out0;
wire  [7:0] v$_15_out0;
wire  [7:0] v$_1644_out0;
wire  [7:0] v$_1645_out0;
wire  [7:0] v$_1646_out0;
wire  [7:0] v$_1647_out0;
wire  [7:0] v$_1648_out0;
wire  [7:0] v$_1649_out0;
wire  [7:0] v$_1650_out0;
wire  [7:0] v$_1651_out0;
wire  [7:0] v$_1652_out0;
wire  [7:0] v$_1653_out0;
wire  [7:0] v$_1654_out0;
wire  [7:0] v$_2023_out0;
wire  [7:0] v$_2068_out0;
wire  [7:0] v$_2315_out0;
wire  [7:0] v$_2316_out0;
wire  [7:0] v$_2378_out1;
wire  [7:0] v$_2379_out1;
wire  [7:0] v$_2424_out0;
wire  [7:0] v$_2489_out1;
wire  [7:0] v$_2490_out1;
wire  [7:0] v$_2491_out1;
wire  [7:0] v$_2492_out1;
wire  [7:0] v$_2493_out1;
wire  [7:0] v$_2494_out1;
wire  [7:0] v$_2495_out1;
wire  [7:0] v$_2496_out1;
wire  [7:0] v$_2497_out1;
wire  [7:0] v$_2498_out1;
wire  [7:0] v$_2499_out1;
wire  [7:0] v$_2516_out0;
wire  [7:0] v$_3006_out0;
wire  [7:0] v$_3006_out1;
wire  [7:0] v$_3007_out0;
wire  [7:0] v$_3007_out1;
wire  [7:0] v$_3086_out0;
wire  [7:0] v$_3125_out0;
wire  [7:0] v$_3358_out0;
wire  [7:0] v$_3359_out0;
wire  [7:0] v$_3360_out0;
wire  [7:0] v$_3372_out1;
wire  [7:0] v$_3435_out0;
wire  [7:0] v$_3537_out0;
wire  [7:0] v$_3847_out0;
wire  [7:0] v$_3924_out0;
wire  [7:0] v$_3925_out0;
wire  [7:0] v$_4349_out1;
wire  [7:0] v$_4350_out1;
wire  [7:0] v$_745_out0;
wire  [7:0] v$_746_out0;
wire  [7:0] v$_747_out0;
wire  [8:0] v$A_3704_out0;
wire  [8:0] v$A_3705_out0;
wire  [8:0] v$A_3706_out0;
wire  [8:0] v$A_3707_out0;
wire  [8:0] v$B_3711_out0;
wire  [8:0] v$B_3712_out0;
wire  [8:0] v$B_3713_out0;
wire  [8:0] v$B_3714_out0;
wire  [8:0] v$C10_5296_out0;
wire  [8:0] v$C12_4493_out0;
wire  [8:0] v$C7_4637_out0;
wire  [8:0] v$C9_1514_out0;
wire  [8:0] v$C_3601_out0;
wire  [8:0] v$C_3602_out0;
wire  [8:0] v$C_3603_out0;
wire  [8:0] v$C_3604_out0;
wire  [8:0] v$S0_1259_out0;
wire  [8:0] v$S0_1260_out0;
wire  [8:0] v$S0_1261_out0;
wire  [8:0] v$S0_1262_out0;
wire  [8:0] v$S1_4224_out0;
wire  [8:0] v$S1_4225_out0;
wire  [8:0] v$S1_4226_out0;
wire  [8:0] v$S1_4227_out0;
wire  [8:0] v$SEL16_3804_out0;
wire  [8:0] v$SEL17_1907_out0;
wire  [8:0] v$SEL18_1412_out0;
wire  [8:0] v$SEL23_4774_out0;
wire  [8:0] v$SEL25_3032_out0;
wire  [8:0] v$SEL27_2724_out0;
wire  [8:0] v$SEL36_2407_out0;
wire  [8:0] v$SEL37_997_out0;
wire  [8:0] v$SEL39_727_out0;
wire  [8:0] v$SEL69_824_out0;
wire  [8:0] v$SEL73_4687_out0;
wire  [8:0] v$SEL75_158_out0;
wire  [8:0] v$X20_4003_out0;
wire  [8:0] v$X8_4348_out0;
wire  [8:0] v$_1016_out0;
wire  [8:0] v$_106_out0;
wire  [8:0] v$_107_out0;
wire  [8:0] v$_1_out0;
wire  [8:0] v$_216_out0;
wire  [8:0] v$_217_out0;
wire  [8:0] v$_218_out0;
wire  [8:0] v$_219_out0;
wire  [8:0] v$_2254_out0;
wire  [8:0] v$_2309_out1;
wire  [8:0] v$_2670_out1;
wire  [8:0] v$_2671_out1;
wire  [8:0] v$_2888_out1;
wire  [8:0] v$_2889_out1;
wire  [8:0] v$_2890_out1;
wire  [8:0] v$_2891_out1;
wire  [8:0] v$_2892_out1;
wire  [8:0] v$_2893_out1;
wire  [8:0] v$_2894_out1;
wire  [8:0] v$_2895_out1;
wire  [8:0] v$_2896_out1;
wire  [8:0] v$_2897_out1;
wire  [8:0] v$_2898_out1;
wire  [8:0] v$_3003_out0;
wire  [8:0] v$_3078_out0;
wire  [8:0] v$_3864_out0;
wire  [8:0] v$_3865_out0;
wire  [8:0] v$_3866_out0;
wire  [8:0] v$_3867_out0;
wire  [8:0] v$_4016_out0;
wire  [8:0] v$_4320_out0;
wire  [8:0] v$_4766_out0;
wire  [8:0] v$_5048_out1;
wire  [8:0] v$_5049_out1;
wire  [8:0] v$_861_out0;
wire  [9:0] v$A_3568_out0;
wire  [9:0] v$A_3569_out0;
wire  [9:0] v$A_3570_out0;
wire  [9:0] v$A_3571_out0;
wire  [9:0] v$B_3840_out0;
wire  [9:0] v$B_3841_out0;
wire  [9:0] v$B_3842_out0;
wire  [9:0] v$B_3843_out0;
wire  [9:0] v$C10_43_out0;
wire  [9:0] v$C12_3681_out0;
wire  [9:0] v$C12_45_out0;
wire  [9:0] v$C4_268_out0;
wire  [9:0] v$C7_311_out0;
wire  [9:0] v$C9_3863_out0;
wire  [9:0] v$C_4517_out0;
wire  [9:0] v$C_4518_out0;
wire  [9:0] v$C_4519_out0;
wire  [9:0] v$C_4520_out0;
wire  [9:0] v$FRACA_1548_out0;
wire  [9:0] v$FRACA_1732_out0;
wire  [9:0] v$FRACB_3484_out0;
wire  [9:0] v$FRACB_3827_out0;
wire  [9:0] v$MUX7_1172_out0;
wire  [9:0] v$NEWFRAC_3836_out0;
wire  [9:0] v$NEWFRAC_608_out0;
wire  [9:0] v$ROUNDEDBITS_4566_out0;
wire  [9:0] v$S1_4205_out0;
wire  [9:0] v$S1_4206_out0;
wire  [9:0] v$S1_4207_out0;
wire  [9:0] v$S1_4208_out0;
wire  [9:0] v$S2_4315_out0;
wire  [9:0] v$S2_4316_out0;
wire  [9:0] v$S2_4317_out0;
wire  [9:0] v$S2_4318_out0;
wire  [9:0] v$SEL1_2457_out0;
wire  [9:0] v$SEL1_2795_out0;
wire  [9:0] v$SEL2_2921_out0;
wire  [9:0] v$SEL2_970_out0;
wire  [9:0] v$SEL31_5225_out0;
wire  [9:0] v$SEL38_465_out0;
wire  [9:0] v$SEL3_3116_out0;
wire  [9:0] v$SEL3_351_out0;
wire  [9:0] v$SEL41_2794_out0;
wire  [9:0] v$SEL43_1228_out0;
wire  [9:0] v$SEL45_173_out0;
wire  [9:0] v$SEL46_5180_out0;
wire  [9:0] v$SEL4_4503_out0;
wire  [9:0] v$SEL83_2369_out0;
wire  [9:0] v$SEL85_3247_out0;
wire  [9:0] v$SEL86_2965_out0;
wire  [9:0] v$X10_2362_out0;
wire  [9:0] v$X17_1251_out0;
wire  [9:0] v$_1145_out1;
wire  [9:0] v$_1265_out1;
wire  [9:0] v$_1266_out1;
wire  [9:0] v$_1267_out1;
wire  [9:0] v$_1268_out1;
wire  [9:0] v$_1269_out1;
wire  [9:0] v$_1270_out1;
wire  [9:0] v$_1271_out1;
wire  [9:0] v$_1272_out1;
wire  [9:0] v$_1273_out1;
wire  [9:0] v$_1274_out1;
wire  [9:0] v$_1275_out1;
wire  [9:0] v$_1290_out0;
wire  [9:0] v$_1291_out0;
wire  [9:0] v$_1361_out0;
wire  [9:0] v$_1825_out0;
wire  [9:0] v$_1927_out0;
wire  [9:0] v$_2500_out0;
wire  [9:0] v$_3038_out0;
wire  [9:0] v$_3039_out0;
wire  [9:0] v$_3040_out0;
wire  [9:0] v$_3041_out0;
wire  [9:0] v$_3590_out0;
wire  [9:0] v$_3608_out0;
wire  [9:0] v$_3609_out0;
wire  [9:0] v$_3610_out0;
wire  [9:0] v$_3611_out0;
wire  [9:0] v$_3807_out0;
wire  [9:0] v$_3916_out0;
wire  [9:0] v$_4319_out0;
wire  [9:0] v$_4443_out0;
wire  [9:0] v$_4578_out0;
wire  [9:0] v$_4723_out1;
wire  [9:0] v$_4724_out1;
wire  [9:0] v$_4820_out1;
wire  [9:0] v$_4821_out1;
wire  [9:0] v$_4938_out0;
wire  [9:0] v$_691_out0;
wire v$0_1011_out0;
wire v$0_1730_out0;
wire v$0_4363_out0;
wire v$0_4364_out0;
wire v$0_4365_out0;
wire v$0_4489_out0;
wire v$10_170_out0;
wire v$10_1774_out0;
wire v$10_4288_out0;
wire v$10_548_out0;
wire v$10_549_out0;
wire v$11_1205_out0;
wire v$11_4305_out0;
wire v$11_4306_out0;
wire v$11_5022_out0;
wire v$12_2636_out0;
wire v$12_2738_out0;
wire v$12_3049_out0;
wire v$12_5202_out0;
wire v$12_5203_out0;
wire v$13_1171_out0;
wire v$13_3103_out0;
wire v$13_935_out0;
wire v$14_1168_out0;
wire v$14_2190_out0;
wire v$14_4529_out0;
wire v$15_287_out0;
wire v$15_2_out0;
wire v$15_4218_out0;
wire v$16_1807_out0;
wire v$16_2631_out0;
wire v$17_364_out0;
wire v$17_4021_out0;
wire v$18_146_out0;
wire v$18_4283_out0;
wire v$19_240_out0;
wire v$19_506_out0;
wire v$1_1838_out0;
wire v$1_3427_out0;
wire v$1_3428_out0;
wire v$1_3429_out0;
wire v$1_4568_out0;
wire v$1_4806_out0;
wire v$1_4807_out0;
wire v$1_5101_out0;
wire v$20_3698_out0;
wire v$20_3805_out0;
wire v$2_1286_out0;
wire v$2_1456_out0;
wire v$2_1783_out0;
wire v$2_1784_out0;
wire v$2_2917_out0;
wire v$2_2918_out0;
wire v$2_2919_out0;
wire v$2_3042_out0;
wire v$3_2559_out0;
wire v$3_2560_out0;
wire v$3_4626_out0;
wire v$3_4627_out0;
wire v$3_4628_out0;
wire v$3_490_out0;
wire v$3_5238_out0;
wire v$3_875_out0;
wire v$4_1200_out0;
wire v$4_1201_out0;
wire v$4_1202_out0;
wire v$4_2368_out0;
wire v$4_718_out0;
wire v$4_92_out0;
wire v$5_2475_out0;
wire v$5_4083_out0;
wire v$5_4084_out0;
wire v$5_4219_out0;
wire v$5_4220_out0;
wire v$5_4221_out0;
wire v$5_4614_out0;
wire v$5_720_out0;
wire v$6_1563_out0;
wire v$6_324_out0;
wire v$6_3495_out0;
wire v$6_3496_out0;
wire v$6_3497_out0;
wire v$6_4279_out0;
wire v$6_4280_out0;
wire v$6_577_out0;
wire v$7_1058_out0;
wire v$7_1310_out0;
wire v$7_1771_out0;
wire v$7_2174_out0;
wire v$7_2175_out0;
wire v$7_4107_out0;
wire v$7_4108_out0;
wire v$7_4951_out0;
wire v$7_4952_out0;
wire v$7_4953_out0;
wire v$8_1388_out0;
wire v$8_1389_out0;
wire v$8_1684_out0;
wire v$8_1972_out0;
wire v$8_1973_out0;
wire v$8_3011_out0;
wire v$8_401_out0;
wire v$9_2615_out0;
wire v$9_2616_out0;
wire v$9_2870_out0;
wire v$9_3255_out0;
wire v$9_784_out0;
wire v$A0_3432_out0;
wire v$A0_550_out0;
wire v$A0_551_out0;
wire v$A0_552_out0;
wire v$A0_553_out0;
wire v$A0_913_out0;
wire v$A0_914_out0;
wire v$A0_915_out0;
wire v$A0_916_out0;
wire v$A10_3265_out0;
wire v$A10_3265_out1;
wire v$A10_3266_out0;
wire v$A10_3266_out1;
wire v$A10_3267_out0;
wire v$A10_3267_out1;
wire v$A10_3268_out0;
wire v$A10_3268_out1;
wire v$A1_1023_out0;
wire v$A1_1023_out1;
wire v$A1_1123_out1;
wire v$A1_1124_out1;
wire v$A1_1299_out0;
wire v$A1_1299_out1;
wire v$A1_1300_out0;
wire v$A1_1300_out1;
wire v$A1_1301_out0;
wire v$A1_1301_out1;
wire v$A1_1302_out0;
wire v$A1_1302_out1;
wire v$A1_1910_out1;
wire v$A1_2039_out1;
wire v$A1_2125_out1;
wire v$A1_2126_out1;
wire v$A1_2427_out1;
wire v$A1_2902_out1;
wire v$A1_2903_out1;
wire v$A1_304_out0;
wire v$A1_331_out1;
wire v$A1_332_out1;
wire v$A1_3679_out1;
wire v$A1_3715_out0;
wire v$A1_3715_out1;
wire v$A1_3716_out0;
wire v$A1_3716_out1;
wire v$A1_3717_out0;
wire v$A1_3717_out1;
wire v$A1_3718_out0;
wire v$A1_3718_out1;
wire v$A1_3820_out0;
wire v$A1_3821_out0;
wire v$A1_3822_out0;
wire v$A1_3823_out0;
wire v$A1_4358_out1;
wire v$A1_5395_out1;
wire v$A1_731_out0;
wire v$A1_732_out0;
wire v$A1_733_out0;
wire v$A1_734_out0;
wire v$A1_794_out1;
wire v$A2_2130_out0;
wire v$A2_2602_out0;
wire v$A2_2602_out1;
wire v$A2_2603_out0;
wire v$A2_2603_out1;
wire v$A2_2604_out0;
wire v$A2_2604_out1;
wire v$A2_2605_out0;
wire v$A2_2605_out1;
wire v$A2_2728_out0;
wire v$A2_2729_out0;
wire v$A2_2730_out0;
wire v$A2_2731_out0;
wire v$A2_312_out0;
wire v$A2_313_out0;
wire v$A2_314_out0;
wire v$A2_315_out0;
wire v$A2_3190_out0;
wire v$A2_3190_out1;
wire v$A2_4328_out0;
wire v$A2_4328_out1;
wire v$A2_4329_out0;
wire v$A2_4329_out1;
wire v$A2_4330_out0;
wire v$A2_4330_out1;
wire v$A2_4331_out0;
wire v$A2_4331_out1;
wire v$A2_4445_out1;
wire v$A2_528_out1;
wire v$A3_1052_out0;
wire v$A3_1053_out0;
wire v$A3_1054_out0;
wire v$A3_1055_out0;
wire v$A3_2871_out0;
wire v$A3_2871_out1;
wire v$A3_2872_out0;
wire v$A3_2872_out1;
wire v$A3_2873_out0;
wire v$A3_2873_out1;
wire v$A3_2874_out0;
wire v$A3_2874_out1;
wire v$A3_368_out0;
wire v$A3_369_out0;
wire v$A3_370_out0;
wire v$A3_371_out0;
wire v$A3_3731_out0;
wire v$A3_3731_out1;
wire v$A3_491_out0;
wire v$A3_5326_out0;
wire v$A3_5326_out1;
wire v$A3_5327_out0;
wire v$A3_5327_out1;
wire v$A3_5328_out0;
wire v$A3_5328_out1;
wire v$A3_5329_out0;
wire v$A3_5329_out1;
wire v$A4_2220_out0;
wire v$A4_2221_out0;
wire v$A4_2222_out0;
wire v$A4_2223_out0;
wire v$A4_2442_out0;
wire v$A4_2443_out0;
wire v$A4_2444_out0;
wire v$A4_2445_out0;
wire v$A4_3034_out0;
wire v$A4_342_out0;
wire v$A4_342_out1;
wire v$A4_343_out0;
wire v$A4_343_out1;
wire v$A4_344_out0;
wire v$A4_344_out1;
wire v$A4_345_out0;
wire v$A4_345_out1;
wire v$A4_519_out0;
wire v$A4_519_out1;
wire v$A4_520_out0;
wire v$A4_520_out1;
wire v$A4_521_out0;
wire v$A4_521_out1;
wire v$A4_522_out0;
wire v$A4_522_out1;
wire v$A4_541_out0;
wire v$A4_541_out1;
wire v$A5_1759_out0;
wire v$A5_1759_out1;
wire v$A5_2706_out0;
wire v$A5_4639_out0;
wire v$A5_4639_out1;
wire v$A5_4640_out0;
wire v$A5_4640_out1;
wire v$A5_4641_out0;
wire v$A5_4641_out1;
wire v$A5_4642_out0;
wire v$A5_4642_out1;
wire v$A5_4738_out0;
wire v$A5_4739_out0;
wire v$A5_4740_out0;
wire v$A5_4741_out0;
wire v$A5_5011_out0;
wire v$A5_5011_out1;
wire v$A5_5012_out0;
wire v$A5_5012_out1;
wire v$A5_5013_out0;
wire v$A5_5013_out1;
wire v$A5_5014_out0;
wire v$A5_5014_out1;
wire v$A5_50_out0;
wire v$A5_51_out0;
wire v$A5_52_out0;
wire v$A5_53_out0;
wire v$A6_1090_out0;
wire v$A6_1090_out1;
wire v$A6_1091_out0;
wire v$A6_1091_out1;
wire v$A6_1092_out0;
wire v$A6_1092_out1;
wire v$A6_1093_out0;
wire v$A6_1093_out1;
wire v$A6_1656_out0;
wire v$A6_1656_out1;
wire v$A6_1657_out0;
wire v$A6_1657_out1;
wire v$A6_1658_out0;
wire v$A6_1658_out1;
wire v$A6_1659_out0;
wire v$A6_1659_out1;
wire v$A6_2072_out0;
wire v$A6_209_out0;
wire v$A6_210_out0;
wire v$A6_211_out0;
wire v$A6_212_out0;
wire v$A6_3768_out0;
wire v$A6_3769_out0;
wire v$A6_3770_out0;
wire v$A6_3771_out0;
wire v$A6_4050_out0;
wire v$A6_4050_out1;
wire v$A7_1862_out0;
wire v$A7_1862_out1;
wire v$A7_1863_out0;
wire v$A7_1863_out1;
wire v$A7_1864_out0;
wire v$A7_1864_out1;
wire v$A7_1865_out0;
wire v$A7_1865_out1;
wire v$A7_3668_out0;
wire v$A7_3668_out1;
wire v$A7_3669_out0;
wire v$A7_3669_out1;
wire v$A7_3670_out0;
wire v$A7_3670_out1;
wire v$A7_3671_out0;
wire v$A7_3671_out1;
wire v$A7_3868_out0;
wire v$A7_3868_out1;
wire v$A7_4079_out0;
wire v$A7_4163_out0;
wire v$A7_4164_out0;
wire v$A7_4165_out0;
wire v$A7_4166_out0;
wire v$A7_4559_out0;
wire v$A7_4560_out0;
wire v$A7_4561_out0;
wire v$A7_4562_out0;
wire v$A8_1452_out0;
wire v$A8_1453_out0;
wire v$A8_1454_out0;
wire v$A8_1455_out0;
wire v$A8_1556_out0;
wire v$A8_1557_out0;
wire v$A8_1558_out0;
wire v$A8_1559_out0;
wire v$A8_1628_out0;
wire v$A8_1628_out1;
wire v$A8_1629_out0;
wire v$A8_1629_out1;
wire v$A8_1630_out0;
wire v$A8_1630_out1;
wire v$A8_1631_out0;
wire v$A8_1631_out1;
wire v$A8_3700_out0;
wire v$A8_3700_out1;
wire v$A8_3701_out0;
wire v$A8_3701_out1;
wire v$A8_3702_out0;
wire v$A8_3702_out1;
wire v$A8_3703_out0;
wire v$A8_3703_out1;
wire v$A9_1280_out0;
wire v$A9_1281_out0;
wire v$A9_1282_out0;
wire v$A9_1283_out0;
wire v$A9_1329_out0;
wire v$A9_1329_out1;
wire v$A9_3763_out0;
wire v$A9_3763_out1;
wire v$A9_3764_out0;
wire v$A9_3764_out1;
wire v$A9_3765_out0;
wire v$A9_3765_out1;
wire v$A9_3766_out0;
wire v$A9_3766_out1;
wire v$A9_4399_out0;
wire v$A9_4399_out1;
wire v$A9_4400_out0;
wire v$A9_4400_out1;
wire v$A9_4401_out0;
wire v$A9_4401_out1;
wire v$A9_4402_out0;
wire v$A9_4402_out1;
wire v$ABEQUAL_2065_out0;
wire v$ABEQUAL_341_out0;
wire v$ABIGGER_2412_out0;
wire v$ABIGGER_4745_out0;
wire v$ABIGGER_4757_out0;
wire v$ADC_1287_out0;
wire v$ADC_1288_out0;
wire v$ADC_3104_out0;
wire v$ADC_3105_out0;
wire v$ADDB_3280_out0;
wire v$ADDONEA_1550_out0;
wire v$ADDONEB_2625_out0;
wire v$ADD_3399_out0;
wire v$ADD_3400_out0;
wire v$ADD_4927_out0;
wire v$ADD_4928_out0;
wire v$ADD_497_out0;
wire v$AND_2179_out0;
wire v$AND_2180_out0;
wire v$AND_46_out0;
wire v$AND_47_out0;
wire v$ASIGN_1780_out0;
wire v$ASMALLER_2055_out0;
wire v$ASMALLER_4525_out0;
wire v$ASMALLER_4819_out0;
wire v$A_2182_out0;
wire v$A_2566_out0;
wire v$A_3523_out0;
wire v$A_4970_out0;
wire v$A_4971_out0;
wire v$A_4972_out0;
wire v$A_4973_out0;
wire v$A_4974_out0;
wire v$A_4975_out0;
wire v$A_4976_out0;
wire v$A_4977_out0;
wire v$A_4978_out0;
wire v$A_4979_out0;
wire v$A_4980_out0;
wire v$A_4981_out0;
wire v$A_4982_out0;
wire v$A_4983_out0;
wire v$A_4984_out0;
wire v$A_4985_out0;
wire v$A_4986_out0;
wire v$A_4987_out0;
wire v$A_4988_out0;
wire v$A_4989_out0;
wire v$A_4990_out0;
wire v$A_4991_out0;
wire v$A_4992_out0;
wire v$A_4993_out0;
wire v$A_4994_out0;
wire v$A_4995_out0;
wire v$A_4996_out0;
wire v$A_4997_out0;
wire v$A_4998_out0;
wire v$Asmaller_2247_out0;
wire v$B0_4340_out0;
wire v$B0_4341_out0;
wire v$B0_4342_out0;
wire v$B0_4343_out0;
wire v$B0_5313_out0;
wire v$B0_5314_out0;
wire v$B0_5315_out0;
wire v$B0_5316_out0;
wire v$B0_5331_out0;
wire v$B1_1748_out0;
wire v$B1_3235_out0;
wire v$B1_3236_out0;
wire v$B1_3237_out0;
wire v$B1_3238_out0;
wire v$B1_5322_out0;
wire v$B1_5323_out0;
wire v$B1_5324_out0;
wire v$B1_5325_out0;
wire v$B2_2645_out0;
wire v$B2_2646_out0;
wire v$B2_2647_out0;
wire v$B2_2648_out0;
wire v$B2_3532_out0;
wire v$B2_764_out0;
wire v$B2_765_out0;
wire v$B2_766_out0;
wire v$B2_767_out0;
wire v$B3_5122_out0;
wire v$B3_5123_out0;
wire v$B3_5124_out0;
wire v$B3_5125_out0;
wire v$B3_705_out0;
wire v$B3_876_out0;
wire v$B3_877_out0;
wire v$B3_878_out0;
wire v$B3_879_out0;
wire v$B4_1867_out0;
wire v$B4_1868_out0;
wire v$B4_1869_out0;
wire v$B4_1870_out0;
wire v$B4_2249_out0;
wire v$B4_2250_out0;
wire v$B4_2251_out0;
wire v$B4_2252_out0;
wire v$B4_2468_out0;
wire v$B5_2656_out0;
wire v$B5_3027_out0;
wire v$B5_3028_out0;
wire v$B5_3029_out0;
wire v$B5_3030_out0;
wire v$B5_4004_out0;
wire v$B5_4005_out0;
wire v$B5_4006_out0;
wire v$B5_4007_out0;
wire v$B6_2662_out0;
wire v$B6_2663_out0;
wire v$B6_2664_out0;
wire v$B6_2665_out0;
wire v$B6_346_out0;
wire v$B6_4850_out0;
wire v$B6_4851_out0;
wire v$B6_4852_out0;
wire v$B6_4853_out0;
wire v$B7_2160_out0;
wire v$B7_2161_out0;
wire v$B7_2162_out0;
wire v$B7_2163_out0;
wire v$B7_3401_out0;
wire v$B7_3918_out0;
wire v$B7_3919_out0;
wire v$B7_3920_out0;
wire v$B7_3921_out0;
wire v$B8_2201_out0;
wire v$B8_2202_out0;
wire v$B8_2203_out0;
wire v$B8_2204_out0;
wire v$B8_3054_out0;
wire v$B8_3055_out0;
wire v$B8_3056_out0;
wire v$B8_3057_out0;
wire v$B9_1440_out0;
wire v$B9_1441_out0;
wire v$B9_1442_out0;
wire v$B9_1443_out0;
wire v$BIGALUSIGN_1581_out0;
wire v$B_147_out0;
wire v$B_3507_out0;
wire v$B_3508_out0;
wire v$B_3509_out0;
wire v$B_3510_out0;
wire v$B_3511_out0;
wire v$B_3512_out0;
wire v$B_3513_out0;
wire v$B_3514_out0;
wire v$B_3515_out0;
wire v$B_3516_out0;
wire v$B_3517_out0;
wire v$B_3975_out0;
wire v$B_4780_out0;
wire v$B_60_out0;
wire v$B_61_out0;
wire v$B_62_out0;
wire v$B_63_out0;
wire v$B_64_out0;
wire v$B_65_out0;
wire v$B_66_out0;
wire v$B_67_out0;
wire v$B_68_out0;
wire v$B_69_out0;
wire v$B_70_out0;
wire v$B_71_out0;
wire v$B_72_out0;
wire v$B_73_out0;
wire v$B_74_out0;
wire v$B_75_out0;
wire v$B_76_out0;
wire v$B_77_out0;
wire v$B_78_out0;
wire v$B_79_out0;
wire v$B_80_out0;
wire v$B_81_out0;
wire v$B_82_out0;
wire v$B_83_out0;
wire v$B_84_out0;
wire v$B_85_out0;
wire v$B_86_out0;
wire v$B_87_out0;
wire v$B_88_out0;
wire v$C0_1107_out0;
wire v$C0_1108_out0;
wire v$C0_1109_out0;
wire v$C0_1110_out0;
wire v$C0_2686_out0;
wire v$C0_419_out0;
wire v$C0_4802_out0;
wire v$C0_5419_out0;
wire v$C0_5420_out0;
wire v$C0_5421_out0;
wire v$C0_5422_out0;
wire v$C14_3974_out0;
wire v$C14_4932_out0;
wire v$C14_4933_out0;
wire v$C15_3806_out0;
wire v$C19_4917_out0;
wire v$C19_4918_out0;
wire v$C1_1176_out0;
wire v$C1_1177_out0;
wire v$C1_1229_out0;
wire v$C1_1230_out0;
wire v$C1_1360_out0;
wire v$C1_1390_out0;
wire v$C1_1391_out0;
wire v$C1_1392_out0;
wire v$C1_1393_out0;
wire v$C1_2702_out0;
wire v$C1_2789_out0;
wire v$C1_3612_out0;
wire v$C1_3691_out0;
wire v$C1_3692_out0;
wire v$C1_3693_out0;
wire v$C1_3694_out0;
wire v$C1_3797_out0;
wire v$C1_3798_out0;
wire v$C1_4332_out0;
wire v$C1_4333_out0;
wire v$C1_5097_out0;
wire v$C1_5098_out0;
wire v$C1_5356_out0;
wire v$C21_4967_out0;
wire v$C23_979_out0;
wire v$C2_1970_out0;
wire v$C2_197_out0;
wire v$C2_198_out0;
wire v$C2_199_out0;
wire v$C2_200_out0;
wire v$C2_23_out0;
wire v$C2_3074_out0;
wire v$C2_3075_out0;
wire v$C2_3989_out0;
wire v$C2_3990_out0;
wire v$C2_3991_out0;
wire v$C2_3992_out0;
wire v$C2_4034_out0;
wire v$C2_5280_out0;
wire v$C2_620_out0;
wire v$C2_621_out0;
wire v$C32_2090_out0;
wire v$C3_2105_out0;
wire v$C3_27_out0;
wire v$C3_28_out0;
wire v$C3_29_out0;
wire v$C3_30_out0;
wire v$C3_3433_out0;
wire v$C3_3579_out0;
wire v$C3_4001_out0;
wire v$C3_4002_out0;
wire v$C3_4732_out0;
wire v$C3_4733_out0;
wire v$C3_4734_out0;
wire v$C3_4735_out0;
wire v$C4_1000_out0;
wire v$C4_1217_out0;
wire v$C4_1218_out0;
wire v$C4_2185_out0;
wire v$C4_3418_out0;
wire v$C4_3419_out0;
wire v$C4_3420_out0;
wire v$C4_3421_out0;
wire v$C4_4228_out0;
wire v$C4_4229_out0;
wire v$C4_4230_out0;
wire v$C4_4231_out0;
wire v$C4_4252_out0;
wire v$C5_1682_out0;
wire v$C5_3631_out0;
wire v$C5_3632_out0;
wire v$C5_3633_out0;
wire v$C5_3634_out0;
wire v$C5_4291_out0;
wire v$C5_4435_out0;
wire v$C5_4513_out0;
wire v$C5_4629_out0;
wire v$C5_4630_out0;
wire v$C5_4631_out0;
wire v$C5_4632_out0;
wire v$C6_1683_out0;
wire v$C6_2674_out0;
wire v$C6_2675_out0;
wire v$C6_2676_out0;
wire v$C6_2677_out0;
wire v$C6_297_out0;
wire v$C6_5170_out0;
wire v$C6_5171_out0;
wire v$C6_5172_out0;
wire v$C6_5173_out0;
wire v$C6_702_out0;
wire v$C7_2317_out0;
wire v$C7_2318_out0;
wire v$C7_2319_out0;
wire v$C7_2320_out0;
wire v$C7_4222_out0;
wire v$C7_4232_out0;
wire v$C7_4233_out0;
wire v$C7_4234_out0;
wire v$C7_4235_out0;
wire v$C7_5135_out0;
wire v$C8_1437_out0;
wire v$C8_2448_out0;
wire v$C8_2449_out0;
wire v$C8_2450_out0;
wire v$C8_2451_out0;
wire v$C8_4120_out0;
wire v$C8_4923_out0;
wire v$C8_4924_out0;
wire v$C8_4925_out0;
wire v$C8_4926_out0;
wire v$C9_697_out0;
wire v$C9_698_out0;
wire v$C9_699_out0;
wire v$C9_700_out0;
wire v$CIN_3082_out0;
wire v$CIN_3083_out0;
wire v$CMP_1059_out0;
wire v$CMP_1060_out0;
wire v$CMP_3183_out0;
wire v$CMP_3184_out0;
wire v$CONTEXTSAVEN_5332_out0;
wire v$CONTEXTSAVEN_5333_out0;
wire v$CONTROLGRANT1_1378_out0;
wire v$CONTROLGRANT1_1722_out0;
wire v$CONTROLGRANT2_406_out0;
wire v$CONTROLGRANT2_4822_out0;
wire v$CONTROLGRANT_1832_out0;
wire v$CONTROLGRANT_1833_out0;
wire v$CONTROLREQ1_3719_out0;
wire v$CONTROLREQ2_5432_out0;
wire v$COUT_1150_out0;
wire v$COUT_1151_out0;
wire v$COUT_3301_out0;
wire v$COUT_3302_out0;
wire v$COUT_4071_out0;
wire v$CYC1_3443_out0;
wire v$CYC1_3894_out0;
wire v$CYC2_1461_out0;
wire v$CYC2_2652_out0;
wire v$CYC2_333_out0;
wire v$CYC2_674_out0;
wire v$C_1100_out0;
wire v$C_1101_out0;
wire v$C_1132_out0;
wire v$C_1133_out0;
wire v$C_2643_out0;
wire v$C_2644_out0;
wire v$C_638_out0;
wire v$C_639_out0;
wire v$C_640_out0;
wire v$C_641_out0;
wire v$C_642_out0;
wire v$C_643_out0;
wire v$C_644_out0;
wire v$C_645_out0;
wire v$C_646_out0;
wire v$C_647_out0;
wire v$C_648_out0;
wire v$C_649_out0;
wire v$C_650_out0;
wire v$C_651_out0;
wire v$C_652_out0;
wire v$C_653_out0;
wire v$C_654_out0;
wire v$C_655_out0;
wire v$C_656_out0;
wire v$C_657_out0;
wire v$C_658_out0;
wire v$C_659_out0;
wire v$C_660_out0;
wire v$C_661_out0;
wire v$C_662_out0;
wire v$C_663_out0;
wire v$C_664_out0;
wire v$C_665_out0;
wire v$C_666_out0;
wire v$C_903_out0;
wire v$C_904_out0;
wire v$D1_3759_out0;
wire v$D1_3759_out1;
wire v$D1_3759_out2;
wire v$D1_3759_out3;
wire v$D1_3760_out0;
wire v$D1_3760_out1;
wire v$D1_3760_out2;
wire v$D1_3760_out3;
wire v$DETECT1_1926_out0;
wire v$DETECT1_2843_out0;
wire v$DETECT1_4467_out0;
wire v$DETECT1_5247_out0;
wire v$DM1_4074_out0;
wire v$DM1_4074_out1;
wire v$DM1_4075_out0;
wire v$DM1_4075_out1;
wire v$DM2_1095_out0;
wire v$DM2_1095_out1;
wire v$EN_1424_out0;
wire v$EN_1425_out0;
wire v$EN_3825_out0;
wire v$EN_3826_out0;
wire v$EN_4955_out0;
wire v$EN_4956_out0;
wire v$EN_5416_out0;
wire v$EN_5417_out0;
wire v$EQ0_4033_out0;
wire v$EQ10_3887_out0;
wire v$EQ10_4417_out0;
wire v$EQ10_5239_out0;
wire v$EQ11_1119_out0;
wire v$EQ11_3818_out0;
wire v$EQ11_707_out0;
wire v$EQ12_1524_out0;
wire v$EQ12_2481_out0;
wire v$EQ13_5289_out0;
wire v$EQ13_963_out0;
wire v$EQ14_785_out0;
wire v$EQ15_2420_out0;
wire v$EQ15_2421_out0;
wire v$EQ15_4014_out0;
wire v$EQ16_329_out0;
wire v$EQ16_330_out0;
wire v$EQ16_564_out0;
wire v$EQ17_35_out0;
wire v$EQ17_719_out0;
wire v$EQ18_1971_out0;
wire v$EQ18_3008_out0;
wire v$EQ19_4433_out0;
wire v$EQ1_1314_out0;
wire v$EQ1_1315_out0;
wire v$EQ1_1321_out0;
wire v$EQ1_1858_out0;
wire v$EQ1_2628_out0;
wire v$EQ1_2629_out0;
wire v$EQ1_2704_out0;
wire v$EQ1_2759_out0;
wire v$EQ1_3286_out0;
wire v$EQ1_3574_out0;
wire v$EQ1_3645_out0;
wire v$EQ1_3646_out0;
wire v$EQ1_4689_out0;
wire v$EQ1_4690_out0;
wire v$EQ1_4746_out0;
wire v$EQ1_4874_out0;
wire v$EQ1_5213_out0;
wire v$EQ1_5269_out0;
wire v$EQ1_5270_out0;
wire v$EQ1_737_out0;
wire v$EQ1_738_out0;
wire v$EQ20_1460_out0;
wire v$EQ21_4249_out0;
wire v$EQ22_1837_out0;
wire v$EQ24_1543_out0;
wire v$EQ25_1034_out0;
wire v$EQ26_4856_out0;
wire v$EQ2_1471_out0;
wire v$EQ2_2556_out0;
wire v$EQ2_2557_out0;
wire v$EQ2_2691_out0;
wire v$EQ2_3018_out0;
wire v$EQ2_3106_out0;
wire v$EQ2_3619_out0;
wire v$EQ2_4098_out0;
wire v$EQ2_4118_out0;
wire v$EQ2_4119_out0;
wire v$EQ2_5128_out0;
wire v$EQ2_5129_out0;
wire v$EQ2_5208_out0;
wire v$EQ2_5209_out0;
wire v$EQ3_1928_out0;
wire v$EQ3_1929_out0;
wire v$EQ3_3053_out0;
wire v$EQ3_3281_out0;
wire v$EQ3_3655_out0;
wire v$EQ3_4099_out0;
wire v$EQ3_4100_out0;
wire v$EQ3_415_out0;
wire v$EQ3_4403_out0;
wire v$EQ3_4404_out0;
wire v$EQ3_4431_out0;
wire v$EQ3_5255_out0;
wire v$EQ4_2879_out0;
wire v$EQ4_2880_out0;
wire v$EQ4_3762_out0;
wire v$EQ4_3781_out0;
wire v$EQ4_4213_out0;
wire v$EQ4_5183_out0;
wire v$EQ4_5388_out0;
wire v$EQ5_1611_out0;
wire v$EQ5_1612_out0;
wire v$EQ5_1712_out0;
wire v$EQ5_3264_out0;
wire v$EQ5_3791_out0;
wire v$EQ5_3879_out0;
wire v$EQ5_4729_out0;
wire v$EQ5_694_out0;
wire v$EQ6_1208_out0;
wire v$EQ6_3613_out0;
wire v$EQ6_3614_out0;
wire v$EQ6_3801_out0;
wire v$EQ6_4710_out0;
wire v$EQ6_4783_out0;
wire v$EQ6_612_out0;
wire v$EQ7_1017_out0;
wire v$EQ7_1762_out0;
wire v$EQ7_2205_out0;
wire v$EQ7_2953_out0;
wire v$EQ7_379_out0;
wire v$EQ7_425_out0;
wire v$EQ7_426_out0;
wire v$EQ8_3303_out0;
wire v$EQ8_3440_out0;
wire v$EQ8_3736_out0;
wire v$EQ8_3737_out0;
wire v$EQ8_504_out0;
wire v$EQ8_5195_out0;
wire v$EQ9_2253_out0;
wire v$EQ9_2267_out0;
wire v$EQ9_2487_out0;
wire v$EQ9_901_out0;
wire v$EQUAL_5338_out0;
wire v$EQUAL_5339_out0;
wire v$EQ_1529_out0;
wire v$EQ_1530_out0;
wire v$EQ_2306_out0;
wire v$EQ_2307_out0;
wire v$EQ_3344_out0;
wire v$EQ_3345_out0;
wire v$EQ_923_out0;
wire v$EQ_924_out0;
wire v$EXCEPTION_1020_out0;
wire v$EXCEPTION_1252_out0;
wire v$EXCEPTION_1402_out0;
wire v$EXCEPTION_1689_out0;
wire v$EXCEPTION_321_out0;
wire v$EXCEPTION_5275_out0;
wire v$EXCEPTION_855_out0;
wire v$EXEC1_201_out0;
wire v$EXEC1_202_out0;
wire v$EXEC1_2363_out0;
wire v$EXEC1_2364_out0;
wire v$EXEC1_2956_out0;
wire v$EXEC1_2957_out0;
wire v$EXEC1_3460_out0;
wire v$EXEC1_3461_out0;
wire v$EXEC1_3733_out0;
wire v$EXEC1_3734_out0;
wire v$EXEC1_3981_out0;
wire v$EXEC1_3982_out0;
wire v$EXEC1_4080_out0;
wire v$EXEC1_4081_out0;
wire v$EXEC2_1668_out0;
wire v$EXEC2_1669_out0;
wire v$EXEC2_1703_out0;
wire v$EXEC2_1704_out0;
wire v$EXEC2_2224_out0;
wire v$EXEC2_2225_out0;
wire v$EXEC2_2321_out0;
wire v$EXEC2_2322_out0;
wire v$EXEC2_3776_out0;
wire v$EXEC2_3777_out0;
wire v$EXEC2_4061_out0;
wire v$EXEC2_4062_out0;
wire v$EXEC2_4334_out0;
wire v$EXEC2_4335_out0;
wire v$EXEC2_4383_out0;
wire v$EXEC2_4384_out0;
wire v$EXEC2_5106_out0;
wire v$EXEC2_5107_out0;
wire v$EXEC2_543_out0;
wire v$EXEC2_544_out0;
wire v$EXEC2_562_out0;
wire v$EXEC2_563_out0;
wire v$EXPOBIGGER_2482_out0;
wire v$EXPOBIGGER_2483_out0;
wire v$EXPONOCHANGE_278_out0;
wire v$F1_5396_out0;
wire v$F2_288_out0;
wire v$FETCH_2291_out0;
wire v$FETCH_2292_out0;
wire v$FETCH_2877_out0;
wire v$FETCH_2878_out0;
wire v$FETCH_3722_out0;
wire v$FETCH_3723_out0;
wire v$FETCH_921_out0;
wire v$FETCH_922_out0;
wire v$FRACTIONINTA_348_out0;
wire v$FRACTIONINTA_631_out0;
wire v$FRACTIONINTB_1578_out0;
wire v$FRACTIONINTB_3004_out0;
wire v$G0_1974_out0;
wire v$G0_1975_out0;
wire v$G0_1976_out0;
wire v$G0_1977_out0;
wire v$G0_1978_out0;
wire v$G0_1979_out0;
wire v$G0_1980_out0;
wire v$G0_1981_out0;
wire v$G0_1982_out0;
wire v$G0_1983_out0;
wire v$G0_1984_out0;
wire v$G0_1985_out0;
wire v$G0_1986_out0;
wire v$G0_1987_out0;
wire v$G0_1988_out0;
wire v$G0_1989_out0;
wire v$G0_1990_out0;
wire v$G0_1991_out0;
wire v$G0_1992_out0;
wire v$G0_1993_out0;
wire v$G0_1994_out0;
wire v$G0_1995_out0;
wire v$G0_1996_out0;
wire v$G0_1997_out0;
wire v$G0_1998_out0;
wire v$G0_1999_out0;
wire v$G0_2000_out0;
wire v$G0_2001_out0;
wire v$G0_2002_out0;
wire v$G10_2259_out0;
wire v$G10_2260_out0;
wire v$G10_2910_out0;
wire v$G10_2911_out0;
wire v$G10_3145_out0;
wire v$G10_3146_out0;
wire v$G10_3240_out0;
wire v$G10_3241_out0;
wire v$G10_5141_out0;
wire v$G10_5142_out0;
wire v$G10_59_out0;
wire v$G11_110_out0;
wire v$G11_111_out0;
wire v$G11_1316_out0;
wire v$G11_1317_out0;
wire v$G11_2141_out0;
wire v$G11_2142_out0;
wire v$G11_4253_out0;
wire v$G11_4254_out0;
wire v$G11_4586_out0;
wire v$G11_4587_out0;
wire v$G11_4588_out0;
wire v$G11_4589_out0;
wire v$G11_4590_out0;
wire v$G11_4591_out0;
wire v$G11_4592_out0;
wire v$G11_4593_out0;
wire v$G11_4594_out0;
wire v$G11_4595_out0;
wire v$G11_4596_out0;
wire v$G11_5397_out0;
wire v$G12_2209_out0;
wire v$G12_2210_out0;
wire v$G12_2211_out0;
wire v$G12_2212_out0;
wire v$G12_2213_out0;
wire v$G12_2214_out0;
wire v$G12_2215_out0;
wire v$G12_2216_out0;
wire v$G12_2217_out0;
wire v$G12_2218_out0;
wire v$G12_2219_out0;
wire v$G12_3199_out0;
wire v$G12_3200_out0;
wire v$G12_5211_out0;
wire v$G12_5212_out0;
wire v$G12_5243_out0;
wire v$G12_5244_out0;
wire v$G13_2037_out0;
wire v$G13_2038_out0;
wire v$G13_254_out0;
wire v$G13_326_out0;
wire v$G13_327_out0;
wire v$G14_1860_out0;
wire v$G14_1861_out0;
wire v$G14_2733_out0;
wire v$G14_285_out0;
wire v$G14_286_out0;
wire v$G14_5078_out0;
wire v$G14_5079_out0;
wire v$G14_5080_out0;
wire v$G14_5081_out0;
wire v$G14_5082_out0;
wire v$G14_5083_out0;
wire v$G14_5084_out0;
wire v$G14_5085_out0;
wire v$G14_5086_out0;
wire v$G14_5087_out0;
wire v$G14_5088_out0;
wire v$G15_1113_out0;
wire v$G15_2300_out0;
wire v$G15_2301_out0;
wire v$G15_2567_out0;
wire v$G15_2568_out0;
wire v$G15_2569_out0;
wire v$G15_2570_out0;
wire v$G15_2571_out0;
wire v$G15_2572_out0;
wire v$G15_2573_out0;
wire v$G15_2574_out0;
wire v$G15_2575_out0;
wire v$G15_2576_out0;
wire v$G15_2577_out0;
wire v$G15_4791_out0;
wire v$G16_1803_out0;
wire v$G16_1804_out0;
wire v$G16_2159_out0;
wire v$G16_890_out0;
wire v$G16_891_out0;
wire v$G16_892_out0;
wire v$G16_893_out0;
wire v$G16_894_out0;
wire v$G16_895_out0;
wire v$G16_896_out0;
wire v$G16_897_out0;
wire v$G16_898_out0;
wire v$G16_899_out0;
wire v$G16_900_out0;
wire v$G16_971_out0;
wire v$G17_1082_out0;
wire v$G17_1083_out0;
wire v$G18_2013_out0;
wire v$G18_2014_out0;
wire v$G19_786_out0;
wire v$G19_787_out0;
wire v$G1_1085_out0;
wire v$G1_1086_out0;
wire v$G1_1184_out0;
wire v$G1_1185_out0;
wire v$G1_1258_out0;
wire v$G1_1886_out0;
wire v$G1_1887_out0;
wire v$G1_1924_out0;
wire v$G1_1925_out0;
wire v$G1_2517_out0;
wire v$G1_2518_out0;
wire v$G1_2519_out0;
wire v$G1_2520_out0;
wire v$G1_2521_out0;
wire v$G1_2522_out0;
wire v$G1_2523_out0;
wire v$G1_2524_out0;
wire v$G1_2525_out0;
wire v$G1_2526_out0;
wire v$G1_2527_out0;
wire v$G1_2528_out0;
wire v$G1_2529_out0;
wire v$G1_2530_out0;
wire v$G1_2531_out0;
wire v$G1_2532_out0;
wire v$G1_2533_out0;
wire v$G1_2534_out0;
wire v$G1_2535_out0;
wire v$G1_2536_out0;
wire v$G1_2537_out0;
wire v$G1_2538_out0;
wire v$G1_2539_out0;
wire v$G1_2540_out0;
wire v$G1_2541_out0;
wire v$G1_2542_out0;
wire v$G1_2543_out0;
wire v$G1_2544_out0;
wire v$G1_2545_out0;
wire v$G1_2775_out0;
wire v$G1_2776_out0;
wire v$G1_2777_out0;
wire v$G1_2778_out0;
wire v$G1_2779_out0;
wire v$G1_2780_out0;
wire v$G1_2781_out0;
wire v$G1_2782_out0;
wire v$G1_2783_out0;
wire v$G1_2784_out0;
wire v$G1_2785_out0;
wire v$G1_2937_out0;
wire v$G1_3684_out0;
wire v$G1_373_out0;
wire v$G1_3741_out0;
wire v$G1_3742_out0;
wire v$G1_3963_out0;
wire v$G1_3964_out0;
wire v$G1_3986_out0;
wire v$G1_4094_out0;
wire v$G1_5051_out0;
wire v$G1_554_out0;
wire v$G1_555_out0;
wire v$G1_695_out0;
wire v$G1_706_out0;
wire v$G1_795_out0;
wire v$G1_909_out0;
wire v$G1_910_out0;
wire v$G1_983_out0;
wire v$G1_984_out0;
wire v$G20_318_out0;
wire v$G20_319_out0;
wire v$G21_1800_out0;
wire v$G21_1801_out0;
wire v$G22_3336_out0;
wire v$G22_3337_out0;
wire v$G23_1484_out0;
wire v$G23_1485_out0;
wire v$G24_2700_out0;
wire v$G24_2701_out0;
wire v$G26_818_out0;
wire v$G26_819_out0;
wire v$G2_1233_out0;
wire v$G2_1242_out0;
wire v$G2_1760_out0;
wire v$G2_1761_out0;
wire v$G2_2236_out0;
wire v$G2_2237_out0;
wire v$G2_2927_out0;
wire v$G2_2928_out0;
wire v$G2_299_out0;
wire v$G2_3352_out0;
wire v$G2_3353_out0;
wire v$G2_3757_out0;
wire v$G2_3758_out0;
wire v$G2_4167_out0;
wire v$G2_4168_out0;
wire v$G2_429_out0;
wire v$G2_430_out0;
wire v$G2_431_out0;
wire v$G2_432_out0;
wire v$G2_433_out0;
wire v$G2_434_out0;
wire v$G2_435_out0;
wire v$G2_436_out0;
wire v$G2_437_out0;
wire v$G2_438_out0;
wire v$G2_439_out0;
wire v$G2_440_out0;
wire v$G2_441_out0;
wire v$G2_442_out0;
wire v$G2_443_out0;
wire v$G2_444_out0;
wire v$G2_445_out0;
wire v$G2_446_out0;
wire v$G2_447_out0;
wire v$G2_448_out0;
wire v$G2_4494_out0;
wire v$G2_449_out0;
wire v$G2_450_out0;
wire v$G2_451_out0;
wire v$G2_452_out0;
wire v$G2_453_out0;
wire v$G2_454_out0;
wire v$G2_455_out0;
wire v$G2_456_out0;
wire v$G2_457_out0;
wire v$G2_4803_out0;
wire v$G2_5045_out0;
wire v$G2_5046_out0;
wire v$G2_518_out0;
wire v$G2_5351_out0;
wire v$G2_5400_out0;
wire v$G2_704_out0;
wire v$G2_721_out0;
wire v$G2_722_out0;
wire v$G2_763_out0;
wire v$G39_1318_out0;
wire v$G39_1319_out0;
wire v$G3_1413_out0;
wire v$G3_1542_out0;
wire v$G3_2173_out0;
wire v$G3_2198_out0;
wire v$G3_2199_out0;
wire v$G3_2338_out0;
wire v$G3_2339_out0;
wire v$G3_2802_out0;
wire v$G3_2803_out0;
wire v$G3_2804_out0;
wire v$G3_2805_out0;
wire v$G3_2806_out0;
wire v$G3_2807_out0;
wire v$G3_2808_out0;
wire v$G3_2809_out0;
wire v$G3_2810_out0;
wire v$G3_2811_out0;
wire v$G3_2812_out0;
wire v$G3_2813_out0;
wire v$G3_2814_out0;
wire v$G3_2815_out0;
wire v$G3_2816_out0;
wire v$G3_2817_out0;
wire v$G3_2818_out0;
wire v$G3_2819_out0;
wire v$G3_2820_out0;
wire v$G3_2821_out0;
wire v$G3_2822_out0;
wire v$G3_2823_out0;
wire v$G3_2824_out0;
wire v$G3_2825_out0;
wire v$G3_2826_out0;
wire v$G3_2827_out0;
wire v$G3_2828_out0;
wire v$G3_2829_out0;
wire v$G3_2830_out0;
wire v$G3_2968_out0;
wire v$G3_3253_out0;
wire v$G3_3254_out0;
wire v$G3_3356_out0;
wire v$G3_3357_out0;
wire v$G3_3467_out0;
wire v$G3_3808_out0;
wire v$G3_4378_out0;
wire v$G3_4379_out0;
wire v$G3_4849_out0;
wire v$G3_5000_out0;
wire v$G3_5001_out0;
wire v$G3_5002_out0;
wire v$G3_5003_out0;
wire v$G3_5004_out0;
wire v$G3_5005_out0;
wire v$G3_5006_out0;
wire v$G3_5007_out0;
wire v$G3_5008_out0;
wire v$G3_5009_out0;
wire v$G3_5010_out0;
wire v$G3_5425_out0;
wire v$G3_6_out0;
wire v$G3_7_out0;
wire v$G40_2289_out0;
wire v$G40_2290_out0;
wire v$G41_1466_out0;
wire v$G41_1467_out0;
wire v$G41_1468_out0;
wire v$G42_2707_out0;
wire v$G42_2708_out0;
wire v$G43_2433_out0;
wire v$G43_2434_out0;
wire v$G43_2435_out0;
wire v$G44_3209_out0;
wire v$G44_3210_out0;
wire v$G44_3211_out0;
wire v$G45_2791_out0;
wire v$G45_2792_out0;
wire v$G45_2793_out0;
wire v$G46_559_out0;
wire v$G46_560_out0;
wire v$G46_561_out0;
wire v$G47_4373_out0;
wire v$G47_4374_out0;
wire v$G47_4375_out0;
wire v$G48_2725_out0;
wire v$G48_2726_out0;
wire v$G48_2727_out0;
wire v$G49_3412_out0;
wire v$G49_3413_out0;
wire v$G49_3414_out0;
wire v$G4_1102_out0;
wire v$G4_1330_out0;
wire v$G4_1331_out0;
wire v$G4_1332_out0;
wire v$G4_1333_out0;
wire v$G4_1334_out0;
wire v$G4_1335_out0;
wire v$G4_1336_out0;
wire v$G4_1337_out0;
wire v$G4_1338_out0;
wire v$G4_1339_out0;
wire v$G4_1340_out0;
wire v$G4_1341_out0;
wire v$G4_1342_out0;
wire v$G4_1343_out0;
wire v$G4_1344_out0;
wire v$G4_1345_out0;
wire v$G4_1346_out0;
wire v$G4_1347_out0;
wire v$G4_1348_out0;
wire v$G4_1349_out0;
wire v$G4_1350_out0;
wire v$G4_1351_out0;
wire v$G4_1352_out0;
wire v$G4_1353_out0;
wire v$G4_1354_out0;
wire v$G4_1355_out0;
wire v$G4_1356_out0;
wire v$G4_1357_out0;
wire v$G4_1358_out0;
wire v$G4_1418_out0;
wire v$G4_2282_out0;
wire v$G4_2283_out0;
wire v$G4_2999_out0;
wire v$G4_3958_out0;
wire v$G4_4284_out0;
wire v$G4_4285_out0;
wire v$G4_4292_out0;
wire v$G4_4293_out0;
wire v$G4_4294_out0;
wire v$G4_4295_out0;
wire v$G4_4296_out0;
wire v$G4_4297_out0;
wire v$G4_4298_out0;
wire v$G4_4299_out0;
wire v$G4_4300_out0;
wire v$G4_4301_out0;
wire v$G4_4302_out0;
wire v$G4_4501_out0;
wire v$G4_4502_out0;
wire v$G4_4548_out0;
wire v$G4_4549_out0;
wire v$G4_4572_out0;
wire v$G4_4743_out0;
wire v$G4_4744_out0;
wire v$G4_5249_out0;
wire v$G4_5336_out0;
wire v$G4_597_out0;
wire v$G4_615_out0;
wire v$G50_246_out0;
wire v$G50_247_out0;
wire v$G50_248_out0;
wire v$G51_3595_out0;
wire v$G51_3596_out0;
wire v$G51_3597_out0;
wire v$G52_301_out0;
wire v$G52_302_out0;
wire v$G52_303_out0;
wire v$G53_2295_out0;
wire v$G53_2296_out0;
wire v$G53_2297_out0;
wire v$G54_2008_out0;
wire v$G54_2009_out0;
wire v$G54_2010_out0;
wire v$G55_3407_out0;
wire v$G55_3408_out0;
wire v$G55_3409_out0;
wire v$G56_2854_out0;
wire v$G56_2855_out0;
wire v$G56_2856_out0;
wire v$G57_4883_out0;
wire v$G57_4884_out0;
wire v$G57_4885_out0;
wire v$G58_4583_out0;
wire v$G58_4584_out0;
wire v$G58_4585_out0;
wire v$G5_1623_out0;
wire v$G5_1876_out0;
wire v$G5_1877_out0;
wire v$G5_2063_out0;
wire v$G5_2945_out0;
wire v$G5_3298_out0;
wire v$G5_3518_out0;
wire v$G5_3519_out0;
wire v$G5_3849_out0;
wire v$G5_3850_out0;
wire v$G5_3851_out0;
wire v$G5_3852_out0;
wire v$G5_3853_out0;
wire v$G5_3854_out0;
wire v$G5_3855_out0;
wire v$G5_3856_out0;
wire v$G5_3857_out0;
wire v$G5_3858_out0;
wire v$G5_3859_out0;
wire v$G5_4111_out0;
wire v$G5_4434_out0;
wire v$G5_5029_out0;
wire v$G5_5030_out0;
wire v$G5_5319_out0;
wire v$G5_5320_out0;
wire v$G5_5359_out0;
wire v$G5_5360_out0;
wire v$G5_5361_out0;
wire v$G5_5362_out0;
wire v$G5_5363_out0;
wire v$G5_5364_out0;
wire v$G5_5365_out0;
wire v$G5_5366_out0;
wire v$G5_5367_out0;
wire v$G5_5368_out0;
wire v$G5_5369_out0;
wire v$G5_5370_out0;
wire v$G5_5371_out0;
wire v$G5_5372_out0;
wire v$G5_5373_out0;
wire v$G5_5374_out0;
wire v$G5_5375_out0;
wire v$G5_5376_out0;
wire v$G5_5377_out0;
wire v$G5_5378_out0;
wire v$G5_5379_out0;
wire v$G5_5380_out0;
wire v$G5_5381_out0;
wire v$G5_5382_out0;
wire v$G5_5383_out0;
wire v$G5_5384_out0;
wire v$G5_5385_out0;
wire v$G5_5386_out0;
wire v$G5_5387_out0;
wire v$G5_729_out0;
wire v$G5_730_out0;
wire v$G60_5426_out0;
wire v$G60_5427_out0;
wire v$G60_5428_out0;
wire v$G61_3941_out0;
wire v$G61_3942_out0;
wire v$G61_3943_out0;
wire v$G62_4941_out0;
wire v$G62_4942_out0;
wire v$G62_4943_out0;
wire v$G63_821_out0;
wire v$G63_822_out0;
wire v$G63_823_out0;
wire v$G64_2688_out0;
wire v$G64_2689_out0;
wire v$G64_2690_out0;
wire v$G65_130_out0;
wire v$G65_131_out0;
wire v$G66_557_out0;
wire v$G66_558_out0;
wire v$G6_1567_out0;
wire v$G6_1568_out0;
wire v$G6_2012_out0;
wire v$G6_2973_out0;
wire v$G6_2974_out0;
wire v$G6_3165_out0;
wire v$G6_3166_out0;
wire v$G6_3167_out0;
wire v$G6_3168_out0;
wire v$G6_3169_out0;
wire v$G6_3170_out0;
wire v$G6_3171_out0;
wire v$G6_3172_out0;
wire v$G6_3173_out0;
wire v$G6_3174_out0;
wire v$G6_3175_out0;
wire v$G6_3367_out0;
wire v$G6_3368_out0;
wire v$G6_3552_out0;
wire v$G6_410_out0;
wire v$G6_411_out0;
wire v$G6_4354_out0;
wire v$G6_4355_out0;
wire v$G6_4376_out0;
wire v$G6_4510_out0;
wire v$G6_4511_out0;
wire v$G6_4830_out0;
wire v$G7_1633_out0;
wire v$G7_1634_out0;
wire v$G7_1635_out0;
wire v$G7_1636_out0;
wire v$G7_1637_out0;
wire v$G7_1638_out0;
wire v$G7_1639_out0;
wire v$G7_1640_out0;
wire v$G7_1641_out0;
wire v$G7_1642_out0;
wire v$G7_1643_out0;
wire v$G7_2835_out0;
wire v$G7_2850_out0;
wire v$G7_3779_out0;
wire v$G7_3780_out0;
wire v$G7_4011_out0;
wire v$G7_4012_out0;
wire v$G7_4776_out0;
wire v$G7_4777_out0;
wire v$G7_5039_out0;
wire v$G7_5040_out0;
wire v$G7_5185_out0;
wire v$G7_5186_out0;
wire v$G8_1121_out0;
wire v$G8_1122_out0;
wire v$G8_1311_out0;
wire v$G8_2419_out0;
wire v$G8_2713_out0;
wire v$G8_2714_out0;
wire v$G8_2899_out0;
wire v$G8_2900_out0;
wire v$G8_4101_out0;
wire v$G8_4102_out0;
wire v$G8_4860_out0;
wire v$G8_4861_out0;
wire v$G9_1426_out0;
wire v$G9_1427_out0;
wire v$G9_3695_out0;
wire v$G9_3696_out0;
wire v$G9_4109_out0;
wire v$G9_4110_out0;
wire v$G9_4580_out0;
wire v$G9_4581_out0;
wire v$G9_5174_out0;
wire v$G9_5175_out0;
wire v$G9_567_out0;
wire v$G9_91_out0;
wire v$IJUMP_1376_out0;
wire v$IJUMP_1377_out0;
wire v$INFINITY16_2098_out0;
wire v$INFINITY2_4485_out0;
wire v$INFINITYA_2940_out0;
wire v$INFINITYB_1096_out0;
wire v$INFINITYB_1517_out0;
wire v$INFINITY_1025_out0;
wire v$INFINITY_2028_out0;
wire v$INFINITY_231_out0;
wire v$INFINITY_4150_out0;
wire v$INTERRUPT1_2431_out0;
wire v$INTERRUPT2_4761_out0;
wire v$INTERRUPT_3178_out0;
wire v$INTERRUPT_3179_out0;
wire v$INTERRUPT_4487_out0;
wire v$INTERRUPT_4488_out0;
wire v$INTERRUPT_93_out0;
wire v$INTERRUPT_94_out0;
wire v$INT_3598_out0;
wire v$IR15_2859_out0;
wire v$IR15_2860_out0;
wire v$IR15_322_out0;
wire v$IR15_323_out0;
wire v$JEQN_2145_out0;
wire v$JEQN_2146_out0;
wire v$JEQN_3047_out0;
wire v$JEQN_3048_out0;
wire v$JMIN_234_out0;
wire v$JMIN_235_out0;
wire v$JMIN_2697_out0;
wire v$JMIN_2698_out0;
wire v$JMPN_1036_out0;
wire v$JMPN_1037_out0;
wire v$JMPN_1855_out0;
wire v$JMPN_1856_out0;
wire v$JMP_2029_out0;
wire v$JMP_2030_out0;
wire v$LOAD_1490_out0;
wire v$LOAD_2672_out0;
wire v$L_1597_out0;
wire v$L_1598_out0;
wire v$MI_1295_out0;
wire v$MI_1296_out0;
wire v$MI_1823_out0;
wire v$MI_1824_out0;
wire v$MI_3185_out0;
wire v$MI_3186_out0;
wire v$MI_4847_out0;
wire v$MI_4848_out0;
wire v$MOV_1952_out0;
wire v$MOV_1953_out0;
wire v$MOV_3738_out0;
wire v$MOV_3739_out0;
wire v$MSB_1458_out0;
wire v$MSB_4908_out0;
wire v$MULTB_3304_out0;
wire v$MULTISHIFT_2679_out0;
wire v$MULT_1828_out0;
wire v$MULT_49_out0;
wire v$MULT_991_out0;
wire v$MUX15_4624_out0;
wire v$MUX15_4625_out0;
wire v$MUX16_3996_out0;
wire v$MUX16_3997_out0;
wire v$MUX17_1733_out0;
wire v$MUX17_1734_out0;
wire v$MUX18_5025_out0;
wire v$MUX18_5026_out0;
wire v$MUX1_3538_out0;
wire v$MUX1_3730_out0;
wire v$MUX2_155_out0;
wire v$MUX2_1594_out0;
wire v$MUX2_1595_out0;
wire v$MUX2_2396_out0;
wire v$MUX2_2397_out0;
wire v$MUX2_3319_out0;
wire v$MUX2_3320_out0;
wire v$MUX2_3778_out0;
wire v$MUX2_4845_out0;
wire v$MUX2_4846_out0;
wire v$MUX2_843_out0;
wire v$MUX3_2226_out0;
wire v$MUX3_3424_out0;
wire v$MUX3_3425_out0;
wire v$MUX3_4659_out0;
wire v$MUX3_4660_out0;
wire v$MUX3_4875_out0;
wire v$MUX3_4876_out0;
wire v$MUX3_693_out0;
wire v$MUX4_3084_out0;
wire v$MUX4_3085_out0;
wire v$MUX5_2340_out0;
wire v$MUX5_2341_out0;
wire v$MUX6_2954_out0;
wire v$MUX6_2955_out0;
wire v$MUX6_572_out0;
wire v$MUX7_2479_out0;
wire v$MUX7_2480_out0;
wire v$MUX8_2410_out0;
wire v$MUX8_2411_out0;
wire v$MUX8_2951_out0;
wire v$MUX8_2952_out0;
wire v$NA_1199_out0;
wire v$NA_4715_out0;
wire v$NA_4716_out0;
wire v$NB_547_out0;
wire v$NEGATIVEMODE_394_out0;
wire v$NEGATIVEMODE_5050_out0;
wire v$NEWSIGN_3096_out0;
wire v$NONVALID_1544_out0;
wire v$NONVALID_3848_out0;
wire v$NONVALID_424_out0;
wire v$NOR_3258_out0;
wire v$NOR_3259_out0;
wire v$NOTUSE10_2286_out0;
wire v$NOTUSE11_3709_out0;
wire v$NOTUSE12_947_out0;
wire v$NOTUSE13_3468_out0;
wire v$NOTUSE1_4377_out0;
wire v$NOTUSE4_1839_out0;
wire v$NOTUSE5_3950_out0;
wire v$NOTUSE6_2721_out0;
wire v$NOTUSE7_2361_out0;
wire v$NOTUSE8_5140_out0;
wire v$NOTUSE9_5190_out0;
wire v$NOTUSED_4919_out0;
wire v$NOTUSED_4920_out0;
wire v$NOTUSEMSB_4611_out0;
wire v$NOTUSE_2079_out0;
wire v$NOTUSE_3678_out0;
wire v$NQ0_5_out0;
wire v$OVERFLOW0_5258_out0;
wire v$OVERFLOW1_4085_out0;
wire v$OVERFLOW_2597_out0;
wire v$OVERFLOW_2773_out0;
wire v$OVERFLOW_2960_out0;
wire v$PRIORITY1_2673_out0;
wire v$PRIORITY2_4698_out0;
wire v$PRIORITYCODE_501_out0;
wire v$PRIORITYCODE_502_out0;
wire v$PRIORITYSAME_5355_out0;
wire v$PRIORITY_2626_out0;
wire v$PRIORITY_2627_out0;
wire v$P_905_out0;
wire v$P_906_out0;
wire v$Q$_2632_out0;
wire v$Q0_356_out0;
wire v$Q_1495_out0;
wire v$RAMWEN_3187_out0;
wire v$RAMWEN_3188_out0;
wire v$READREQ_2930_out0;
wire v$READREQ_2931_out0;
wire v$READREQ_5066_out0;
wire v$READREQ_5067_out0;
wire v$READVALID_178_out0;
wire v$READVALID_179_out0;
wire v$READVALID_2915_out0;
wire v$READVALID_2916_out0;
wire v$RET_2021_out0;
wire v$RET_2022_out0;
wire v$RET_2085_out0;
wire v$RET_2086_out0;
wire v$RET_2207_out0;
wire v$RET_2208_out0;
wire v$RET_2238_out0;
wire v$RET_2239_out0;
wire v$RET_3361_out0;
wire v$RET_3362_out0;
wire v$RET_4161_out0;
wire v$RET_4162_out0;
wire v$RET_4312_out0;
wire v$RET_4313_out0;
wire v$RET_622_out0;
wire v$RET_623_out0;
wire v$RET_677_out0;
wire v$RET_678_out0;
wire v$RIGHTSHIFT_4693_out0;
wire v$RREQUEST_3720_out0;
wire v$RREQUEST_3721_out0;
wire v$S00_1128_out0;
wire v$S00_1129_out0;
wire v$S00_1130_out0;
wire v$S00_1131_out0;
wire v$S00_2884_out0;
wire v$S00_4439_out0;
wire v$S00_4440_out0;
wire v$S00_4441_out0;
wire v$S00_4442_out0;
wire v$S01_1061_out0;
wire v$S01_1062_out0;
wire v$S01_1063_out0;
wire v$S01_1064_out0;
wire v$S01_191_out0;
wire v$S01_192_out0;
wire v$S01_193_out0;
wire v$S01_194_out0;
wire v$S01_5221_out0;
wire v$S02_1072_out0;
wire v$S02_1073_out0;
wire v$S02_1074_out0;
wire v$S02_1075_out0;
wire v$S02_1187_out0;
wire v$S02_3390_out0;
wire v$S02_3391_out0;
wire v$S02_3392_out0;
wire v$S02_3393_out0;
wire v$S03_2844_out0;
wire v$S03_2845_out0;
wire v$S03_2846_out0;
wire v$S03_2847_out0;
wire v$S03_3014_out0;
wire v$S03_3015_out0;
wire v$S03_3016_out0;
wire v$S03_3017_out0;
wire v$S03_4045_out0;
wire v$S04_2278_out0;
wire v$S04_2279_out0;
wire v$S04_2280_out0;
wire v$S04_2281_out0;
wire v$S04_4731_out0;
wire v$S04_927_out0;
wire v$S04_928_out0;
wire v$S04_929_out0;
wire v$S04_930_out0;
wire v$S05_2988_out0;
wire v$S05_2989_out0;
wire v$S05_2990_out0;
wire v$S05_2991_out0;
wire v$S05_3458_out0;
wire v$S05_4886_out0;
wire v$S05_4887_out0;
wire v$S05_4888_out0;
wire v$S05_4889_out0;
wire v$S06_3111_out0;
wire v$S06_3112_out0;
wire v$S06_3113_out0;
wire v$S06_3114_out0;
wire v$S06_3373_out0;
wire v$S06_4367_out0;
wire v$S06_4368_out0;
wire v$S06_4369_out0;
wire v$S06_4370_out0;
wire v$S07_1254_out0;
wire v$S07_1255_out0;
wire v$S07_1256_out0;
wire v$S07_1257_out0;
wire v$S07_5042_out0;
wire v$S07_886_out0;
wire v$S07_887_out0;
wire v$S07_888_out0;
wire v$S07_889_out0;
wire v$S08_1589_out0;
wire v$S08_1590_out0;
wire v$S08_1591_out0;
wire v$S08_1592_out0;
wire v$S08_5271_out0;
wire v$S08_5272_out0;
wire v$S08_5273_out0;
wire v$S08_5274_out0;
wire v$S09_1936_out0;
wire v$S09_1937_out0;
wire v$S09_1938_out0;
wire v$S09_1939_out0;
wire v$S10_3263_out0;
wire v$S10_3471_out0;
wire v$S10_3472_out0;
wire v$S10_3473_out0;
wire v$S10_3474_out0;
wire v$S10_938_out0;
wire v$S10_939_out0;
wire v$S10_940_out0;
wire v$S10_941_out0;
wire v$S11_2561_out0;
wire v$S11_2562_out0;
wire v$S11_2563_out0;
wire v$S11_2564_out0;
wire v$S11_3140_out0;
wire v$S11_3141_out0;
wire v$S11_3142_out0;
wire v$S11_3143_out0;
wire v$S11_3803_out0;
wire v$S12_100_out0;
wire v$S12_101_out0;
wire v$S12_102_out0;
wire v$S12_103_out0;
wire v$S12_4495_out0;
wire v$S12_4798_out0;
wire v$S12_4799_out0;
wire v$S12_4800_out0;
wire v$S12_4801_out0;
wire v$S13_1157_out0;
wire v$S13_3436_out0;
wire v$S13_3437_out0;
wire v$S13_3438_out0;
wire v$S13_3439_out0;
wire v$S13_851_out0;
wire v$S13_852_out0;
wire v$S13_853_out0;
wire v$S13_854_out0;
wire v$S14_3379_out0;
wire v$S14_3380_out0;
wire v$S14_3381_out0;
wire v$S14_3382_out0;
wire v$S14_667_out0;
wire v$S14_668_out0;
wire v$S14_669_out0;
wire v$S14_670_out0;
wire v$S14_753_out0;
wire v$S15_3216_out0;
wire v$S15_3217_out0;
wire v$S15_3218_out0;
wire v$S15_3219_out0;
wire v$S15_458_out0;
wire v$S15_459_out0;
wire v$S15_460_out0;
wire v$S15_461_out0;
wire v$S15_542_out0;
wire v$S16_3242_out0;
wire v$S16_4694_out0;
wire v$S16_4695_out0;
wire v$S16_4696_out0;
wire v$S16_4697_out0;
wire v$S16_4891_out0;
wire v$S16_4892_out0;
wire v$S16_4893_out0;
wire v$S16_4894_out0;
wire v$S17_2861_out0;
wire v$S17_2862_out0;
wire v$S17_2863_out0;
wire v$S17_2864_out0;
wire v$S17_4090_out0;
wire v$S17_4091_out0;
wire v$S17_4092_out0;
wire v$S17_4093_out0;
wire v$S17_4121_out0;
wire v$S18_1961_out0;
wire v$S18_1962_out0;
wire v$S18_1963_out0;
wire v$S18_1964_out0;
wire v$S18_2436_out0;
wire v$S18_2437_out0;
wire v$S18_2438_out0;
wire v$S18_2439_out0;
wire v$S19_568_out0;
wire v$S19_569_out0;
wire v$S19_570_out0;
wire v$S19_571_out0;
wire v$SBC_2040_out0;
wire v$SBC_2041_out0;
wire v$SBC_4704_out0;
wire v$SBC_4705_out0;
wire v$SEL10_1158_out0;
wire v$SEL10_1159_out0;
wire v$SEL10_1160_out0;
wire v$SEL10_1161_out0;
wire v$SEL10_3410_out0;
wire v$SEL10_4314_out0;
wire v$SEL10_4864_out0;
wire v$SEL10_4865_out0;
wire v$SEL10_4866_out0;
wire v$SEL10_4867_out0;
wire v$SEL11_1602_out0;
wire v$SEL11_2549_out0;
wire v$SEL11_2550_out0;
wire v$SEL11_2551_out0;
wire v$SEL11_2552_out0;
wire v$SEL11_2553_out0;
wire v$SEL11_3134_out0;
wire v$SEL11_3135_out0;
wire v$SEL11_3136_out0;
wire v$SEL11_3137_out0;
wire v$SEL11_3875_out0;
wire v$SEL12_1173_out0;
wire v$SEL12_1174_out0;
wire v$SEL12_2081_out0;
wire v$SEL12_2082_out0;
wire v$SEL12_2083_out0;
wire v$SEL12_2084_out0;
wire v$SEL12_2598_out0;
wire v$SEL12_3895_out0;
wire v$SEL12_4139_out0;
wire v$SEL12_4140_out0;
wire v$SEL12_4141_out0;
wire v$SEL12_4142_out0;
wire v$SEL13_2981_out0;
wire v$SEL13_2982_out0;
wire v$SEL13_2983_out0;
wire v$SEL13_2984_out0;
wire v$SEL13_3455_out0;
wire v$SEL13_3456_out0;
wire v$SEL13_3457_out0;
wire v$SEL13_3869_out0;
wire v$SEL13_3870_out0;
wire v$SEL13_3871_out0;
wire v$SEL13_3872_out0;
wire v$SEL13_3911_out0;
wire v$SEL13_4643_out0;
wire v$SEL14_1153_out0;
wire v$SEL14_1154_out0;
wire v$SEL14_1155_out0;
wire v$SEL14_1491_out0;
wire v$SEL14_1492_out0;
wire v$SEL14_1493_out0;
wire v$SEL14_1494_out0;
wire v$SEL14_4787_out0;
wire v$SEL14_5214_out0;
wire v$SEL14_5215_out0;
wire v$SEL14_5216_out0;
wire v$SEL14_5217_out0;
wire v$SEL15_1363_out0;
wire v$SEL15_1364_out0;
wire v$SEL15_1365_out0;
wire v$SEL15_1366_out0;
wire v$SEL15_467_out0;
wire v$SEL15_468_out0;
wire v$SEL15_469_out0;
wire v$SEL15_4950_out0;
wire v$SEL15_496_out0;
wire v$SEL15_830_out0;
wire v$SEL15_831_out0;
wire v$SEL15_832_out0;
wire v$SEL15_833_out0;
wire v$SEL16_1170_out0;
wire v$SEL16_1895_out0;
wire v$SEL16_1896_out0;
wire v$SEL16_1897_out0;
wire v$SEL16_1898_out0;
wire v$SEL16_2266_out0;
wire v$SEL16_3937_out0;
wire v$SEL16_3938_out0;
wire v$SEL16_3939_out0;
wire v$SEL16_3940_out0;
wire v$SEL16_4038_out0;
wire v$SEL16_4039_out0;
wire v$SEL16_4040_out0;
wire v$SEL17_3824_out0;
wire v$SEL17_3944_out0;
wire v$SEL17_3945_out0;
wire v$SEL17_3946_out0;
wire v$SEL17_4471_out0;
wire v$SEL17_4472_out0;
wire v$SEL17_4473_out0;
wire v$SEL17_4474_out0;
wire v$SEL17_992_out0;
wire v$SEL17_993_out0;
wire v$SEL17_994_out0;
wire v$SEL17_995_out0;
wire v$SEL18_2406_out0;
wire v$SEL18_24_out0;
wire v$SEL18_25_out0;
wire v$SEL18_26_out0;
wire v$SEL18_3444_out0;
wire v$SEL18_3449_out0;
wire v$SEL18_3450_out0;
wire v$SEL18_3451_out0;
wire v$SEL18_3452_out0;
wire v$SEL18_4245_out0;
wire v$SEL18_4246_out0;
wire v$SEL18_4247_out0;
wire v$SEL18_4248_out0;
wire v$SEL19_1071_out0;
wire v$SEL19_1486_out0;
wire v$SEL19_1487_out0;
wire v$SEL19_1488_out0;
wire v$SEL19_1489_out0;
wire v$SEL19_1532_out0;
wire v$SEL19_1533_out0;
wire v$SEL19_1534_out0;
wire v$SEL19_1535_out0;
wire v$SEL19_3244_out0;
wire v$SEL19_4778_out0;
wire v$SEL1_1279_out0;
wire v$SEL1_2413_out0;
wire v$SEL1_2548_out0;
wire v$SEL1_3201_out0;
wire v$SEL1_3202_out0;
wire v$SEL1_3203_out0;
wire v$SEL1_3204_out0;
wire v$SEL1_3305_out0;
wire v$SEL1_3306_out0;
wire v$SEL1_3307_out0;
wire v$SEL1_3308_out0;
wire v$SEL1_3332_out0;
wire v$SEL1_4138_out0;
wire v$SEL1_4767_out0;
wire v$SEL1_4768_out0;
wire v$SEL1_4771_out0;
wire v$SEL1_4808_out0;
wire v$SEL1_4854_out0;
wire v$SEL1_744_out0;
wire v$SEL20_1841_out0;
wire v$SEL20_1842_out0;
wire v$SEL20_1843_out0;
wire v$SEL20_1844_out0;
wire v$SEL20_2270_out0;
wire v$SEL20_2271_out0;
wire v$SEL20_2272_out0;
wire v$SEL20_4543_out0;
wire v$SEL20_4544_out0;
wire v$SEL20_4545_out0;
wire v$SEL20_4546_out0;
wire v$SEL20_848_out0;
wire v$SEL21_2091_out0;
wire v$SEL21_2092_out0;
wire v$SEL21_2093_out0;
wire v$SEL21_2848_out0;
wire v$SEL21_4308_out0;
wire v$SEL21_4309_out0;
wire v$SEL21_4310_out0;
wire v$SEL21_4311_out0;
wire v$SEL21_754_out0;
wire v$SEL21_755_out0;
wire v$SEL21_756_out0;
wire v$SEL21_757_out0;
wire v$SEL21_969_out0;
wire v$SEL22_1249_out0;
wire v$SEL22_2743_out0;
wire v$SEL22_2922_out0;
wire v$SEL22_2923_out0;
wire v$SEL22_2924_out0;
wire v$SEL22_2925_out0;
wire v$SEL22_514_out0;
wire v$SEL22_958_out0;
wire v$SEL22_959_out0;
wire v$SEL22_960_out0;
wire v$SEL22_961_out0;
wire v$SEL23_3951_out0;
wire v$SEL23_3968_out0;
wire v$SEL23_3969_out0;
wire v$SEL23_3970_out0;
wire v$SEL23_3971_out0;
wire v$SEL23_584_out0;
wire v$SEL23_585_out0;
wire v$SEL23_586_out0;
wire v$SEL23_587_out0;
wire v$SEL23_9_out0;
wire v$SEL24_1407_out0;
wire v$SEL24_1408_out0;
wire v$SEL24_1409_out0;
wire v$SEL24_1410_out0;
wire v$SEL24_1791_out0;
wire v$SEL24_1792_out0;
wire v$SEL24_1793_out0;
wire v$SEL24_1794_out0;
wire v$SEL24_1834_out0;
wire v$SEL24_2372_out0;
wire v$SEL24_3660_out0;
wire v$SEL24_4859_out0;
wire v$SEL25_1731_out0;
wire v$SEL25_402_out0;
wire v$SEL25_4211_out0;
wire v$SEL25_4655_out0;
wire v$SEL25_4656_out0;
wire v$SEL25_4657_out0;
wire v$SEL25_4658_out0;
wire v$SEL25_4719_out0;
wire v$SEL25_4720_out0;
wire v$SEL25_4721_out0;
wire v$SEL25_4722_out0;
wire v$SEL26_1706_out0;
wire v$SEL26_1707_out0;
wire v$SEL26_1708_out0;
wire v$SEL26_1709_out0;
wire v$SEL26_1763_out0;
wire v$SEL26_1764_out0;
wire v$SEL26_1765_out0;
wire v$SEL26_1766_out0;
wire v$SEL26_3130_out0;
wire v$SEL26_3328_out0;
wire v$SEL26_466_out0;
wire v$SEL26_529_out0;
wire v$SEL27_2607_out0;
wire v$SEL27_2608_out0;
wire v$SEL27_2609_out0;
wire v$SEL27_2610_out0;
wire v$SEL27_3260_out0;
wire v$SEL27_412_out0;
wire v$SEL27_917_out0;
wire v$SEL27_918_out0;
wire v$SEL27_919_out0;
wire v$SEL27_920_out0;
wire v$SEL28_143_out0;
wire v$SEL28_3406_out0;
wire v$SEL28_4554_out0;
wire v$SEL28_4555_out0;
wire v$SEL28_4556_out0;
wire v$SEL28_4557_out0;
wire v$SEL29_4444_out0;
wire v$SEL29_4456_out0;
wire v$SEL29_96_out0;
wire v$SEL29_97_out0;
wire v$SEL29_98_out0;
wire v$SEL29_99_out0;
wire v$SEL2_1112_out0;
wire v$SEL2_1234_out0;
wire v$SEL2_1235_out0;
wire v$SEL2_2432_out0;
wire v$SEL2_3384_out0;
wire v$SEL2_3922_out0;
wire v$SEL2_3962_out0;
wire v$SEL2_4366_out0;
wire v$SEL2_4934_out0;
wire v$SEL2_5056_out0;
wire v$SEL2_5204_out0;
wire v$SEL2_5321_out0;
wire v$SEL2_603_out0;
wire v$SEL2_604_out0;
wire v$SEL2_605_out0;
wire v$SEL2_606_out0;
wire v$SEL2_739_out0;
wire v$SEL2_740_out0;
wire v$SEL2_741_out0;
wire v$SEL2_742_out0;
wire v$SEL30_1539_out0;
wire v$SEL30_1613_out0;
wire v$SEL30_1614_out0;
wire v$SEL30_1615_out0;
wire v$SEL30_1616_out0;
wire v$SEL30_2716_out0;
wire v$SEL31_4563_out0;
wire v$SEL32_36_out0;
wire v$SEL32_696_out0;
wire v$SEL33_1035_out0;
wire v$SEL33_1822_out0;
wire v$SEL34_2547_out0;
wire v$SEL35_1547_out0;
wire v$SEL36_3144_out0;
wire v$SEL37_2633_out0;
wire v$SEL38_4463_out0;
wire v$SEL3_1276_out0;
wire v$SEL3_1362_out0;
wire v$SEL3_1482_out0;
wire v$SEL3_1662_out0;
wire v$SEL3_1663_out0;
wire v$SEL3_1664_out0;
wire v$SEL3_1665_out0;
wire v$SEL3_1892_out0;
wire v$SEL3_3088_out0;
wire v$SEL3_357_out0;
wire v$SEL3_358_out0;
wire v$SEL3_359_out0;
wire v$SEL3_360_out0;
wire v$SEL3_4260_out0;
wire v$SEL3_4770_out0;
wire v$SEL3_5279_out0;
wire v$SEL40_4711_out0;
wire v$SEL42_2134_out0;
wire v$SEL42_3888_out0;
wire v$SEL43_1956_out0;
wire v$SEL44_2612_out0;
wire v$SEL46_1049_out0;
wire v$SEL47_1719_out0;
wire v$SEL48_3948_out0;
wire v$SEL49_2881_out0;
wire v$SEL4_2184_out0;
wire v$SEL4_275_out0;
wire v$SEL4_3161_out0;
wire v$SEL4_3162_out0;
wire v$SEL4_3163_out0;
wire v$SEL4_3164_out0;
wire v$SEL4_3355_out0;
wire v$SEL4_38_out0;
wire v$SEL4_39_out0;
wire v$SEL4_40_out0;
wire v$SEL4_41_out0;
wire v$SEL4_464_out0;
wire v$SEL4_5071_out0;
wire v$SEL4_768_out0;
wire v$SEL50_2478_out0;
wire v$SEL50_736_out0;
wire v$SEL53_4486_out0;
wire v$SEL54_4089_out0;
wire v$SEL55_752_out0;
wire v$SEL56_1474_out0;
wire v$SEL57_2938_out0;
wire v$SEL58_4499_out0;
wire v$SEL59_4818_out0;
wire v$SEL5_1596_out0;
wire v$SEL5_1923_out0;
wire v$SEL5_266_out0;
wire v$SEL5_267_out0;
wire v$SEL5_3239_out0;
wire v$SEL5_3697_out0;
wire v$SEL5_3993_out0;
wire v$SEL5_4029_out0;
wire v$SEL5_4030_out0;
wire v$SEL5_4031_out0;
wire v$SEL5_4032_out0;
wire v$SEL5_4146_out0;
wire v$SEL5_4147_out0;
wire v$SEL5_4148_out0;
wire v$SEL5_4149_out0;
wire v$SEL5_4204_out0;
wire v$SEL5_4688_out0;
wire v$SEL5_701_out0;
wire v$SEL63_3931_out0;
wire v$SEL64_2195_out0;
wire v$SEL65_3615_out0;
wire v$SEL66_1553_out0;
wire v$SEL67_815_out0;
wire v$SEL6_1041_out0;
wire v$SEL6_1042_out0;
wire v$SEL6_1043_out0;
wire v$SEL6_1044_out0;
wire v$SEL6_1507_out0;
wire v$SEL6_1508_out0;
wire v$SEL6_1509_out0;
wire v$SEL6_1510_out0;
wire v$SEL6_1560_out0;
wire v$SEL6_1561_out0;
wire v$SEL6_2071_out0;
wire v$SEL6_227_out0;
wire v$SEL6_2599_out0;
wire v$SEL6_3676_out0;
wire v$SEL6_582_out0;
wire v$SEL70_2638_out0;
wire v$SEL71_3374_out0;
wire v$SEL72_215_out0;
wire v$SEL74_1540_out0;
wire v$SEL77_2323_out0;
wire v$SEL78_4371_out0;
wire v$SEL7_105_out0;
wire v$SEL7_1405_out0;
wire v$SEL7_1406_out0;
wire v$SEL7_1847_out0;
wire v$SEL7_1848_out0;
wire v$SEL7_1849_out0;
wire v$SEL7_1850_out0;
wire v$SEL7_2971_out0;
wire v$SEL7_4775_out0;
wire v$SEL7_5191_out0;
wire v$SEL7_5192_out0;
wire v$SEL7_5193_out0;
wire v$SEL7_5194_out0;
wire v$SEL80_1577_out0;
wire v$SEL82_2669_out0;
wire v$SEL84_4290_out0;
wire v$SEL87_244_out0;
wire v$SEL88_4558_out0;
wire v$SEL8_1503_out0;
wire v$SEL8_1504_out0;
wire v$SEL8_1505_out0;
wire v$SEL8_1506_out0;
wire v$SEL8_3411_out0;
wire v$SEL8_352_out0;
wire v$SEL8_355_out0;
wire v$SEL8_4725_out0;
wire v$SEL8_4726_out0;
wire v$SEL8_4727_out0;
wire v$SEL8_4728_out0;
wire v$SEL90_2866_out0;
wire v$SEL9_3315_out0;
wire v$SEL9_3316_out0;
wire v$SEL9_3317_out0;
wire v$SEL9_3318_out0;
wire v$SEL9_3386_out0;
wire v$SEL9_3387_out0;
wire v$SEL9_3388_out0;
wire v$SEL9_3389_out0;
wire v$SEL9_3961_out0;
wire v$SEL9_4261_out0;
wire v$SEL9_507_out0;
wire v$SERIESCONNECT_3100_out0;
wire v$SERIESCONNECT_4605_out0;
wire v$SERIESCONNECT_4606_out0;
wire v$SGNA_3917_out0;
wire v$SGNA_4123_out0;
wire v$SGNBIGALU_3546_out0;
wire v$SGNB_1810_out0;
wire v$SGNB_3492_out0;
wire v$SGNOUT_2961_out0;
wire v$SGN_3620_out0;
wire v$SIGNOPERATION_3729_out0;
wire v$SIGNTOSHIFT_255_out0;
wire v$SIGNTOSHIFT_3033_out0;
wire v$SIGNTOSHIFT_5047_out0;
wire v$SIGN_1005_out0;
wire v$SIGN_5044_out0;
wire v$STALL1_3563_out0;
wire v$STALL2_2936_out0;
wire v$STALL_2382_out0;
wire v$STALL_2383_out0;
wire v$STALL_2680_out0;
wire v$STALL_2681_out0;
wire v$STALL_3987_out0;
wire v$STALL_3988_out0;
wire v$STALL_4418_out0;
wire v$STALL_4419_out0;
wire v$STALL_4480_out0;
wire v$STALL_4481_out0;
wire v$STALL_4645_out0;
wire v$STALL_4646_out0;
wire v$STALL_5064_out0;
wire v$STALL_5065_out0;
wire v$STALL_5393_out0;
wire v$STALL_5394_out0;
wire v$STICKY_1727_out0;
wire v$STORESHADOW_1626_out0;
wire v$STORESHADOW_1627_out0;
wire v$STORESHADOW_1787_out0;
wire v$STORESHADOW_1788_out0;
wire v$STORESHADOW_2370_out0;
wire v$STORESHADOW_2371_out0;
wire v$STORESHADOW_3475_out0;
wire v$STORESHADOW_3476_out0;
wire v$STORESHADOW_3540_out0;
wire v$STORESHADOW_3541_out0;
wire v$STORESHADOW_4961_out0;
wire v$STORESHADOW_4962_out0;
wire v$STORESHADOW_632_out0;
wire v$STORESHADOW_633_out0;
wire v$STORESHADOW_859_out0;
wire v$STORESHADOW_860_out0;
wire v$STP_1717_out0;
wire v$STP_1718_out0;
wire v$STP_2446_out0;
wire v$STP_2447_out0;
wire v$STP_4410_out0;
wire v$STP_4411_out0;
wire v$SUBB_4737_out0;
wire v$SUBTRACTOR_1459_out0;
wire v$SUBTRACTOR_3177_out0;
wire v$SUB_2466_out0;
wire v$SUB_2467_out0;
wire v$SUB_3369_out0;
wire v$SUB_3370_out0;
wire v$SUB_3371_out0;
wire v$SUB_3499_out0;
wire v$SUB_4899_out0;
wire v$SUB_510_out0;
wire v$SUB_5242_out0;
wire v$SWITCH_4096_out0;
wire v$SWITCH_4809_out0;
wire v$S_3348_out0;
wire v$S_3349_out0;
wire v$S_4175_out0;
wire v$S_4176_out0;
wire v$S_4177_out0;
wire v$S_4178_out0;
wire v$S_4179_out0;
wire v$S_4180_out0;
wire v$S_4181_out0;
wire v$S_4182_out0;
wire v$S_4183_out0;
wire v$S_4184_out0;
wire v$S_4185_out0;
wire v$S_4186_out0;
wire v$S_4187_out0;
wire v$S_4188_out0;
wire v$S_4189_out0;
wire v$S_4190_out0;
wire v$S_4191_out0;
wire v$S_4192_out0;
wire v$S_4193_out0;
wire v$S_4194_out0;
wire v$S_4195_out0;
wire v$S_4196_out0;
wire v$S_4197_out0;
wire v$S_4198_out0;
wire v$S_4199_out0;
wire v$S_4200_out0;
wire v$S_4201_out0;
wire v$S_4202_out0;
wire v$S_4203_out0;
wire v$S_4391_out0;
wire v$S_4392_out0;
wire v$TOOSMALL_4217_out0;
wire v$TST_1125_out0;
wire v$TST_1126_out0;
wire v$TST_826_out0;
wire v$TST_827_out0;
wire v$U_1679_out0;
wire v$U_1680_out0;
wire v$U_54_out0;
wire v$U_55_out0;
wire v$WEN3_931_out0;
wire v$WEN3_932_out0;
wire v$WENALU_2753_out0;
wire v$WENALU_2754_out0;
wire v$WENALU_5353_out0;
wire v$WENALU_5354_out0;
wire v$WENLDST_1028_out0;
wire v$WENLDST_1029_out0;
wire v$WENLDST_334_out0;
wire v$WENLDST_335_out0;
wire v$WENRAM_5126_out0;
wire v$WENRAM_5127_out0;
wire v$WREQUEST_508_out0;
wire v$WREQUEST_509_out0;
wire v$WRITECOMPLETE_203_out0;
wire v$WRITECOMPLETE_204_out0;
wire v$WRITECOMPLETE_487_out0;
wire v$WRITECOMPLETE_488_out0;
wire v$WRITEENABLE_3250_out0;
wire v$WRITEENABLE_790_out0;
wire v$WRITEREQ_2132_out0;
wire v$WRITEREQ_2133_out0;
wire v$WRITEREQ_4482_out0;
wire v$WRITEREQ_4483_out0;
wire v$W_1874_out0;
wire v$W_1875_out0;
wire v$X1_1220_out0;
wire v$X1_165_out0;
wire v$X1_4916_out0;
wire v$X5_4793_out0;
wire v$XOR1_679_out0;
wire v$X_1263_out0;
wire v$X_1667_out0;
wire v$X_4262_out0;
wire v$X_4263_out0;
wire v$X_530_out0;
wire v$X_759_out0;
wire v$ZERO14_3688_out0;
wire v$ZERO14_4652_out0;
wire v$ZERO_2473_out0;
wire v$ZERO_778_out0;
wire v$_11_out0;
wire v$_1238_out0;
wire v$_1239_out0;
wire v$_1244_out0;
wire v$_1244_out1;
wire v$_1245_out0;
wire v$_1245_out1;
wire v$_1265_out0;
wire v$_1266_out0;
wire v$_1267_out0;
wire v$_1268_out0;
wire v$_1269_out0;
wire v$_1270_out0;
wire v$_1271_out0;
wire v$_1272_out0;
wire v$_1273_out0;
wire v$_1274_out0;
wire v$_1275_out0;
wire v$_1297_out0;
wire v$_1298_out0;
wire v$_12_out0;
wire v$_1512_out0;
wire v$_1512_out1;
wire v$_1513_out0;
wire v$_1513_out1;
wire v$_1569_out0;
wire v$_1569_out1;
wire v$_1570_out0;
wire v$_1570_out1;
wire v$_1580_out0;
wire v$_1580_out1;
wire v$_1701_out0;
wire v$_1702_out0;
wire v$_1728_out0;
wire v$_1729_out0;
wire v$_1749_out0;
wire v$_1750_out0;
wire v$_180_out0;
wire v$_180_out1;
wire v$_1811_out1;
wire v$_181_out0;
wire v$_181_out1;
wire v$_182_out0;
wire v$_182_out1;
wire v$_183_out0;
wire v$_183_out1;
wire v$_184_out0;
wire v$_184_out1;
wire v$_185_out0;
wire v$_185_out1;
wire v$_186_out0;
wire v$_186_out1;
wire v$_1879_out0;
wire v$_1879_out1;
wire v$_187_out0;
wire v$_187_out1;
wire v$_1880_out0;
wire v$_1880_out1;
wire v$_188_out0;
wire v$_188_out1;
wire v$_189_out0;
wire v$_189_out1;
wire v$_190_out0;
wire v$_190_out1;
wire v$_1927_out1;
wire v$_2006_out1;
wire v$_2111_out0;
wire v$_2112_out0;
wire v$_2113_out0;
wire v$_2114_out0;
wire v$_2115_out0;
wire v$_2116_out0;
wire v$_2117_out0;
wire v$_2118_out0;
wire v$_2119_out0;
wire v$_2120_out0;
wire v$_2121_out0;
wire v$_2148_out0;
wire v$_2149_out0;
wire v$_2150_out0;
wire v$_2151_out0;
wire v$_2152_out0;
wire v$_2153_out0;
wire v$_2154_out0;
wire v$_2155_out0;
wire v$_2156_out0;
wire v$_2157_out0;
wire v$_2158_out0;
wire v$_2186_out0;
wire v$_2186_out1;
wire v$_2187_out0;
wire v$_2187_out1;
wire v$_2196_out0;
wire v$_2197_out0;
wire v$_223_out0;
wire v$_224_out0;
wire v$_2284_out1;
wire v$_2285_out1;
wire v$_2378_out0;
wire v$_2379_out0;
wire v$_242_out0;
wire v$_243_out0;
wire v$_2489_out0;
wire v$_2490_out0;
wire v$_2491_out0;
wire v$_2492_out0;
wire v$_2493_out0;
wire v$_2494_out0;
wire v$_2495_out0;
wire v$_2496_out0;
wire v$_2497_out0;
wire v$_2498_out0;
wire v$_2499_out0;
wire v$_256_out0;
wire v$_257_out0;
wire v$_2586_out0;
wire v$_2587_out0;
wire v$_2588_out0;
wire v$_2589_out0;
wire v$_2590_out0;
wire v$_2591_out0;
wire v$_2592_out0;
wire v$_2593_out0;
wire v$_2594_out0;
wire v$_2595_out0;
wire v$_2596_out0;
wire v$_2623_out0;
wire v$_2624_out0;
wire v$_2670_out0;
wire v$_2671_out0;
wire v$_2687_out0;
wire v$_2717_out0;
wire v$_2718_out0;
wire v$_2747_out0;
wire v$_2748_out0;
wire v$_2760_out0;
wire v$_2761_out0;
wire v$_2865_out1;
wire v$_2888_out0;
wire v$_2889_out0;
wire v$_2890_out0;
wire v$_2891_out0;
wire v$_2892_out0;
wire v$_2893_out0;
wire v$_2894_out0;
wire v$_2895_out0;
wire v$_2896_out0;
wire v$_2897_out0;
wire v$_2898_out0;
wire v$_2949_out0;
wire v$_2950_out0;
wire v$_2987_out1;
wire v$_2993_out0;
wire v$_2994_out0;
wire v$_3126_out0;
wire v$_3127_out0;
wire v$_3191_out0;
wire v$_3191_out1;
wire v$_3192_out0;
wire v$_3192_out1;
wire v$_3335_out0;
wire v$_3365_out1;
wire v$_3464_out0;
wire v$_3464_out1;
wire v$_3534_out1;
wire v$_3535_out1;
wire v$_3667_out0;
wire v$_3745_out0;
wire v$_3746_out0;
wire v$_3747_out0;
wire v$_3748_out0;
wire v$_3749_out0;
wire v$_3750_out0;
wire v$_3751_out0;
wire v$_3752_out0;
wire v$_3753_out0;
wire v$_3754_out0;
wire v$_3755_out0;
wire v$_3772_out0;
wire v$_3773_out0;
wire v$_3782_out0;
wire v$_3782_out1;
wire v$_3783_out0;
wire v$_3783_out1;
wire v$_3832_out1;
wire v$_3833_out1;
wire v$_4077_out0;
wire v$_4078_out0;
wire v$_4236_out0;
wire v$_4236_out1;
wire v$_4237_out0;
wire v$_4237_out1;
wire v$_4250_out0;
wire v$_4251_out0;
wire v$_4344_out0;
wire v$_4344_out1;
wire v$_4345_out0;
wire v$_4345_out1;
wire v$_4349_out0;
wire v$_4350_out0;
wire v$_4420_out0;
wire v$_4421_out0;
wire v$_4422_out0;
wire v$_4423_out0;
wire v$_4424_out0;
wire v$_4425_out0;
wire v$_4426_out0;
wire v$_4427_out0;
wire v$_4428_out0;
wire v$_4429_out0;
wire v$_4430_out0;
wire v$_4457_out0;
wire v$_4457_out1;
wire v$_4458_out0;
wire v$_4458_out1;
wire v$_4633_out0;
wire v$_4634_out0;
wire v$_4723_out0;
wire v$_4724_out0;
wire v$_4748_out0;
wire v$_4804_out0;
wire v$_4805_out0;
wire v$_4820_out0;
wire v$_4821_out0;
wire v$_4832_out0;
wire v$_4833_out0;
wire v$_4834_out0;
wire v$_4835_out0;
wire v$_4836_out0;
wire v$_4837_out0;
wire v$_4838_out0;
wire v$_4839_out0;
wire v$_4840_out0;
wire v$_4841_out0;
wire v$_4842_out0;
wire v$_4906_out0;
wire v$_4907_out0;
wire v$_4931_out0;
wire v$_5027_out0;
wire v$_5028_out0;
wire v$_5048_out0;
wire v$_5049_out0;
wire v$_5062_out1;
wire v$_5063_out1;
wire v$_5096_out0;
wire v$_5099_out0;
wire v$_5100_out0;
wire v$_5143_out0;
wire v$_5143_out1;
wire v$_5144_out0;
wire v$_5144_out1;
wire v$_523_out0;
wire v$_523_out1;
wire v$_524_out0;
wire v$_524_out1;
wire v$_5317_out0;
wire v$_5318_out0;
wire v$_773_out0;
wire v$_774_out0;
wire v$_862_out1;
wire v$_863_out1;
wire v$_880_out0;
wire v$_881_out0;
wire v$comparator_4432_out1;
wire v$interruptatexec2_3984_out0;
wire v$interruptatexec2_3985_out0;
wire v$interruptatexec2_4897_out0;
wire v$interruptatexec2_4898_out0;
wire v$interruptatexec2_5035_out0;
wire v$interruptatexec2_5036_out0;

always @(posedge clk) v$FF4_89_out0 <= v$LOAD_1490_out0;
always @(posedge clk) v$FF1_144_out0 <= v$STALL_2382_out0;
always @(posedge clk) v$FF1_145_out0 <= v$STALL_2383_out0;
always @(posedge clk) v$FF5_271_out0 <= v$READVALID_2915_out0;
always @(posedge clk) v$REG1_374_out0 <= v$G10_3240_out0 ? v$MUX5_2882_out0 : v$REG1_374_out0;
always @(posedge clk) v$REG1_375_out0 <= v$G10_3241_out0 ? v$MUX5_2883_out0 : v$REG1_375_out0;
always @(posedge clk) v$REG3_574_out0 <= v$STORESHADOW_859_out0 ? v$G4_4284_out0 : v$REG3_574_out0;
always @(posedge clk) v$REG3_575_out0 <= v$STORESHADOW_860_out0 ? v$G4_4285_out0 : v$REG3_575_out0;
always @(posedge clk) v$REG2_750_out0 <= v$interruptatexec2_4897_out0 ? v$MUX7_4351_out0 : v$REG2_750_out0;
always @(posedge clk) v$REG2_751_out0 <= v$interruptatexec2_4898_out0 ? v$MUX7_4352_out0 : v$REG2_751_out0;
always @(posedge clk) v$FF1_846_out0 <= v$G4_2999_out0 ? v$G5_3298_out0 : v$FF1_846_out0;
always @(posedge clk) v$REG1_1106_out0 <= v$G8_1311_out0 ? v$MUX2_5187_out0 : v$REG1_1106_out0;
v$RAM3_1304 I1304 (v$RAM3_1304_out0, v$DMADDRESS_1885_out0, v$WRITEDATA_1328_out0, v$WRITEENABLE_790_out0, clk);
always @(posedge clk) v$REG1_1399_out0 <= v$MUX16_3996_out0 ? v$MUX12_152_out0 : v$REG1_1399_out0;
always @(posedge clk) v$REG1_1400_out0 <= v$MUX16_3997_out0 ? v$MUX12_153_out0 : v$REG1_1400_out0;
always @(posedge clk) v$FF1_1575_out0 <= v$_3772_out0;
always @(posedge clk) v$FF1_1576_out0 <= v$_3773_out0;
always @(posedge clk) v$FF1_1618_out0 <= v$_4344_out0;
always @(posedge clk) v$FF1_1619_out0 <= v$_4345_out0;
always @(posedge clk) v$REG4_1772_out0 <= v$CONTEXTSAVEN_5332_out0 ? v$R3_1883_out0 : v$REG4_1772_out0;
always @(posedge clk) v$REG4_1773_out0 <= v$CONTEXTSAVEN_5333_out0 ? v$R3_1884_out0 : v$REG4_1773_out0;
always @(posedge clk) v$FF2_1859_out0 <= v$READVALID_2916_out0;
always @(posedge clk) v$REG2_1904_out0 <= v$STORESHADOW_859_out0 ? v$G1_1886_out0 : v$REG2_1904_out0;
always @(posedge clk) v$REG2_1905_out0 <= v$STORESHADOW_860_out0 ? v$G1_1887_out0 : v$REG2_1905_out0;
always @(posedge clk) v$FF1_2042_out0 <= v$STALL_4645_out0;
always @(posedge clk) v$FF1_2043_out0 <= v$STALL_4646_out0;
always @(posedge clk) v$REG3_2164_out0 <= v$CONTEXTSAVEN_5332_out0 ? v$R2_3009_out0 : v$REG3_2164_out0;
always @(posedge clk) v$REG3_2165_out0 <= v$CONTEXTSAVEN_5333_out0 ? v$R2_3010_out0 : v$REG3_2165_out0;
always @(posedge clk) v$FF1_2233_out0 <= v$Q$_2632_out0;
always @(posedge clk) v$FF2_2554_out0 <= v$STORESHADOW_1626_out0 ? v$FF1_2975_out0 : v$FF2_2554_out0;
always @(posedge clk) v$FF2_2555_out0 <= v$STORESHADOW_1627_out0 ? v$FF1_2976_out0 : v$FF2_2555_out0;
always @(posedge clk) v$REG1_2682_out0 <= v$CONTEXTSAVEN_5332_out0 ? v$R0_1056_out0 : v$REG1_2682_out0;
always @(posedge clk) v$REG1_2683_out0 <= v$CONTEXTSAVEN_5333_out0 ? v$R0_1057_out0 : v$REG1_2683_out0;
always @(posedge clk) v$REG2_2762_out0 <= v$CONTEXTSAVEN_5332_out0 ? v$R1_4338_out0 : v$REG2_2762_out0;
always @(posedge clk) v$REG2_2763_out0 <= v$CONTEXTSAVEN_5333_out0 ? v$R1_4339_out0 : v$REG2_2763_out0;
always @(posedge clk) v$REG3_2962_out0 <= v$MUX18_5025_out0 ? v$MUX14_1674_out0 : v$REG3_2962_out0;
always @(posedge clk) v$REG3_2963_out0 <= v$MUX18_5026_out0 ? v$MUX14_1675_out0 : v$REG3_2963_out0;
always @(posedge clk) v$FF1_2975_out0 <= v$G11_110_out0 ? v$MUX8_2410_out0 : v$FF1_2975_out0;
always @(posedge clk) v$FF1_2976_out0 <= v$G11_111_out0 ? v$MUX8_2411_out0 : v$FF1_2976_out0;
always @(posedge clk) v$REG5_3036_out0 <= v$G10_3145_out0 ? v$RM_3021_out0 : v$REG5_3036_out0;
always @(posedge clk) v$REG5_3037_out0 <= v$G10_3146_out0 ? v$RM_3022_out0 : v$REG5_3037_out0;
always @(posedge clk) v$FF4_3156_out0 <= v$_1569_out1;
always @(posedge clk) v$FF4_3157_out0 <= v$_1570_out1;
always @(posedge clk) v$REG1_3272_out0 <= v$EXEC2_2321_out0 ? v$ALUOUT_1496_out0 : v$REG1_3272_out0;
always @(posedge clk) v$REG1_3273_out0 <= v$EXEC2_2322_out0 ? v$ALUOUT_1497_out0 : v$REG1_3273_out0;
always @(posedge clk) v$FF2_3299_out0 <= v$G14_1860_out0 ? v$INTERRUPT_93_out0 : v$FF2_3299_out0;
always @(posedge clk) v$FF2_3300_out0 <= v$G14_1861_out0 ? v$INTERRUPT_94_out0 : v$FF2_3300_out0;
always @(posedge clk) v$FF2_3403_out0 <= v$MULTB_3304_out0;
always @(posedge clk) v$REG1_3653_out0 <= v$G2_2236_out0 ? v$RAMDOUT_2667_out0 : v$REG1_3653_out0;
always @(posedge clk) v$REG1_3654_out0 <= v$G2_2237_out0 ? v$RAMDOUT_2668_out0 : v$REG1_3654_out0;
v$ROM3_3844 I3844 (v$ROM3_3844_out0, v$PROGRAMADDRESS_4514_out0, clk);
always @(posedge clk) v$FF1_4133_out0 <= v$G4_4743_out0 ? v$INTERRUPT_93_out0 : v$FF1_4133_out0;
always @(posedge clk) v$FF1_4134_out0 <= v$G4_4744_out0 ? v$INTERRUPT_94_out0 : v$FF1_4134_out0;
always @(posedge clk) v$FF2_4169_out0 <= v$_4344_out1;
always @(posedge clk) v$FF2_4170_out0 <= v$_4345_out1;
always @(posedge clk) v$FF2_4405_out0 <= v$_2284_out1;
always @(posedge clk) v$FF2_4406_out0 <= v$_2285_out1;
always @(posedge clk) v$FF3_4436_out0 <= v$_1569_out0;
always @(posedge clk) v$FF3_4437_out0 <= v$_1570_out0;
always @(posedge clk) v$REG0_4539_out0 <= v$MUX15_4624_out0 ? v$MUX11_1403_out0 : v$REG0_4539_out0;
always @(posedge clk) v$REG0_4540_out0 <= v$MUX15_4625_out0 ? v$MUX11_1404_out0 : v$REG0_4540_out0;
always @(posedge clk) v$REG4_4843_out0 <= v$EXEC2_2321_out0 ? v$ALUOUT_1496_out0 : v$REG4_4843_out0;
always @(posedge clk) v$REG4_4844_out0 <= v$EXEC2_2322_out0 ? v$ALUOUT_1497_out0 : v$REG4_4844_out0;
always @(posedge clk) v$REG2_4872_out0 <= v$MUX17_1733_out0 ? v$MUX13_4054_out0 : v$REG2_4872_out0;
always @(posedge clk) v$REG2_4873_out0 <= v$MUX17_1734_out0 ? v$MUX13_4055_out0 : v$REG2_4873_out0;
v$ROM4_4954 I4954 (v$ROM4_4954_out0, v$PROGRAMADDRESS_4515_out0, clk);
always @(posedge clk) v$FF1_5073_out0 <= v$SUBB_4737_out0;
always @(posedge clk) v$REG2_5309_out0 <= v$G16_971_out0 ? v$WDATA_4407_out0 : v$REG2_5309_out0;
assign v$C19_5406_out0 = 5'h9;
assign v$C2_5404_out0 = 16'hffff;
assign v$C2_5403_out0 = 16'hffff;
assign v$C3_5358_out0 = 4'h1;
assign v$C3_5357_out0 = 4'h1;
assign v$C17_5302_out0 = 5'h1;
assign v$C10_5296_out0 = 9'h0;
assign v$C13_5266_out0 = 5'h1;
assign v$C7_5237_out0 = 7'h0;
assign v$C21_5199_out0 = 5'hb;
assign v$C6_5119_out0 = 6'h0;
assign v$C1_5098_out0 = 1'h0;
assign v$C1_5097_out0 = 1'h0;
assign v$C17_5068_out0 = 2'h0;
assign v$C21_4967_out0 = 1'h0;
assign v$C1_4937_out0 = 13'h1fff;
assign v$C14_4933_out0 = 1'h1;
assign v$C14_4932_out0 = 1'h1;
assign v$C19_4918_out0 = 1'h0;
assign v$C19_4917_out0 = 1'h0;
assign v$C28_4909_out0 = 14'h0;
assign v$C3_4882_out0 = 3'h0;
assign v$C20_4877_out0 = 5'h0;
assign v$C6_4824_out0 = 4'h4;
assign v$C6_4823_out0 = 4'h4;
assign v$C0_4802_out0 = 1'h1;
assign v$C1_4681_out0 = 2'h0;
assign v$C22_4676_out0 = 18'h0;
assign v$C5_4673_out0 = 8'h0;
assign v$C7_4637_out0 = 9'h0;
assign v$C3_4571_out0 = 3'h0;
assign v$C2_4547_out0 = 7'h71;
assign v$C5_4513_out0 = 1'h1;
assign v$C12_4493_out0 = 9'h0;
assign v$C3_4484_out0 = 2'h0;
assign v$C5_4465_out0 = 4'h3;
assign v$C5_4464_out0 = 4'h3;
assign v$C2_4460_out0 = 4'h0;
assign v$C2_4459_out0 = 4'h0;
assign v$C5_4435_out0 = 1'h0;
assign v$C11_4416_out0 = 11'h0;
assign v$C1_4333_out0 = 1'h0;
assign v$C1_4332_out0 = 1'h0;
assign v$C1_4327_out0 = 5'h2;
assign v$C9_4326_out0 = 7'h0;
assign v$C5_4307_out0 = 5'h0;
assign v$C30_4304_out0 = 5'h14;
assign v$C5_4291_out0 = 1'h1;
assign v$C5_4278_out0 = 6'h0;
assign v$C15_4273_out0 = 7'h0;
assign v$C7_4222_out0 = 1'h1;
assign v$C5_4214_out0 = 4'h0;
assign v$C21_4143_out0 = 13'h0;
assign v$C8_4137_out0 = 8'h0;
assign v$C24_4122_out0 = 15'h0;
assign v$C8_4120_out0 = 1'h0;
assign v$C8_4082_out0 = 7'h0;
assign v$C29_4076_out0 = 19'h0;
assign v$C2_4034_out0 = 1'h0;
assign v$C1_4010_out0 = 2'h0;
assign v$C1_4009_out0 = 2'h0;
assign v$C3_4002_out0 = 1'h0;
assign v$C3_4001_out0 = 1'h0;
assign v$C14_3974_out0 = 1'h1;
assign v$C11_3973_out0 = 5'h3;
assign v$C6_3912_out0 = 3'h0;
assign v$C18_3898_out0 = 5'h11;
assign v$C15_3897_out0 = 6'h3f;
assign v$C15_3896_out0 = 8'hff;
assign v$C3_3893_out0 = 2'h0;
assign v$C9_3886_out0 = 5'h1;
assign v$C9_3863_out0 = 10'h0;
assign v$C15_3806_out0 = 1'h0;
assign v$C1_3798_out0 = 1'h1;
assign v$C1_3797_out0 = 1'h1;
assign v$C25_3774_out0 = 13'h0;
assign v$C2_3735_out0 = 6'h0;
assign v$C12_3681_out0 = 10'h0;
assign v$C27_3680_out0 = 5'h0;
assign v$C1_3659_out0 = 4'h0;
assign v$C1_3658_out0 = 4'h0;
assign v$C30_3636_out0 = 16'h0;
assign v$C10_3628_out0 = 5'h0;
assign v$C1_3612_out0 = 1'h0;
assign v$C3_3579_out0 = 1'h1;
assign v$C2_3555_out0 = 5'h0;
assign v$C31_3551_out0 = 5'h13;
assign v$C6_3524_out0 = 6'h0;
assign v$C6_3481_out0 = 5'h1f;
assign v$C3_3433_out0 = 1'h0;
assign v$C11_3383_out0 = 4'h0;
assign v$C11_3343_out0 = 4'h9;
assign v$C11_3342_out0 = 4'h9;
assign v$C4_3256_out0 = 5'h8;
assign v$ROR_3252_out0 = 2'h3;
assign v$ROR_3251_out0 = 2'h3;
assign v$C6_3198_out0 = 5'h0;
assign v$C1_3138_out0 = 6'h0;
assign v$C2_3117_out0 = 2'h0;
assign v$C4_3094_out0 = 12'h20;
assign v$C4_3093_out0 = 12'h20;
assign v$C22_3079_out0 = 2'h0;
assign v$C2_3075_out0 = 1'h0;
assign v$C2_3074_out0 = 1'h0;
assign v$C8_3052_out0 = 5'h7;
assign v$C25_3012_out0 = 20'h0;
assign v$C3_3005_out0 = 3'h0;
assign v$C10_2986_out0 = 5'h1;
assign v$C24_2887_out0 = 8'h0;
assign v$C9_2797_out0 = 4'h7;
assign v$C9_2796_out0 = 4'h7;
assign v$C1_2789_out0 = 1'h0;
assign v$C2_2749_out0 = 2'h0;
assign v$C14_2741_out0 = 4'hc;
assign v$C14_2740_out0 = 4'hc;
assign v$C10_2703_out0 = 7'h0;
assign v$C1_2702_out0 = 1'h0;
assign v$C0_2686_out0 = 1'h1;
assign v$C1_2666_out0 = 5'h0;
assign v$C8_2635_out0 = 4'h6;
assign v$C8_2634_out0 = 4'h6;
assign v$C6_2426_out0 = 5'h0;
assign v$C18_2405_out0 = 13'h0;
assign v$C1_2377_out0 = 8'h0;
assign v$C1_2376_out0 = 8'h0;
assign v$C1_2374_out0 = 5'h1f;
assign v$C12_2311_out0 = 4'ha;
assign v$C12_2310_out0 = 4'ha;
assign v$C1_2299_out0 = 4'h0;
assign v$C1_2298_out0 = 4'h0;
assign v$C2_2234_out0 = 5'h1f;
assign v$C1_2206_out0 = 5'h0;
assign v$C5_2191_out0 = 6'h0;
assign v$C4_2185_out0 = 1'h0;
assign v$C15_2147_out0 = 5'hd;
assign v$C32_2090_out0 = 1'h0;
assign v$C4_2077_out0 = 3'h0;
assign v$C7_2066_out0 = 5'h1f;
assign v$C1_2032_out0 = 12'h0;
assign v$C1_2031_out0 = 12'h0;
assign v$C4_2007_out0 = 4'h0;
assign v$C2_1970_out0 = 1'h0;
assign v$C10_1969_out0 = 4'h8;
assign v$C10_1968_out0 = 4'h8;
assign v$C7_1909_out0 = 4'h5;
assign v$C7_1908_out0 = 4'h5;
assign v$C5_1899_out0 = 4'h0;
assign v$C1_1743_out0 = 12'h0;
assign v$C1_1742_out0 = 12'h0;
assign v$C11_1736_out0 = 11'h0;
assign v$C13_1573_out0 = 7'h7f;
assign v$C3_1546_out0 = 16'h0;
assign v$C3_1545_out0 = 16'h0;
assign v$C4_1537_out0 = 8'h0;
assign v$C18_1516_out0 = 2'h0;
assign v$C18_1515_out0 = 3'h0;
assign v$C9_1514_out0 = 9'h0;
assign v$C20_1438_out0 = 5'hc;
assign v$C8_1437_out0 = 1'h0;
assign v$C9_1415_out0 = 5'h1;
assign v$C3_1385_out0 = 5'h5;
assign v$C1_1360_out0 = 1'h0;
assign v$C12_1322_out0 = 5'h4;
assign v$C1_1312_out0 = 11'h7ff;
assign v$C13_1293_out0 = 4'hb;
assign v$C13_1292_out0 = 4'hb;
assign v$C10_1253_out0 = 4'h0;
assign v$C1_1230_out0 = 1'h1;
assign v$C1_1229_out0 = 1'h1;
assign v$C4_1218_out0 = 1'h1;
assign v$C4_1217_out0 = 1'h1;
assign v$C28_1203_out0 = 5'h1;
assign v$C26_1186_out0 = 4'h0;
assign v$C1_1177_out0 = 1'h1;
assign v$C1_1176_out0 = 1'h1;
assign v$C12_1162_out0 = 12'h0;
assign v$C1_1147_out0 = 11'h0;
assign v$C1_1146_out0 = 11'h0;
assign v$C17_1139_out0 = 5'h10;
assign v$C31_1111_out0 = 2'h0;
assign v$C4_1032_out0 = 4'h2;
assign v$C4_1031_out0 = 4'h2;
assign v$C13_1012_out0 = 13'h0;
assign v$C28_1010_out0 = 5'h12;
assign v$C4_1000_out0 = 1'h1;
assign v$C23_979_out0 = 1'h0;
assign v$C1_865_out0 = 16'h0;
assign v$C1_864_out0 = 16'h0;
assign v$C7_825_out0 = 7'h0;
assign v$C26_791_out0 = 17'h0;
assign v$C4_777_out0 = 5'h0;
assign v$C9_758_out0 = 8'h0;
assign v$C2_743_out0 = 13'h0;
assign v$C6_702_out0 = 1'h0;
assign v$C11_671_out0 = 11'h0;
assign v$C4_627_out0 = 3'h0;
assign v$C2_621_out0 = 1'h0;
assign v$C2_620_out0 = 1'h0;
assign v$C8_598_out0 = 8'h0;
assign v$C14_576_out0 = 5'hf;
assign v$C30_536_out0 = 5'h0;
assign v$C16_427_out0 = 5'he;
assign v$C4_396_out0 = 16'hffff;
assign v$C4_395_out0 = 16'hffff;
assign v$C22_372_out0 = 5'ha;
assign v$C8_338_out0 = 2'h0;
assign v$C13_325_out0 = 12'h0;
assign v$C7_311_out0 = 10'h0;
assign v$C6_297_out0 = 1'h0;
assign v$C13_274_out0 = 7'h0;
assign v$C4_268_out0 = 10'h0;
assign v$C7_228_out0 = 6'h0;
assign v$C16_206_out0 = 5'h0;
assign v$C16_205_out0 = 5'h0;
assign v$C12_45_out0 = 10'h0;
assign v$C10_43_out0 = 10'h0;
assign v$C6_34_out0 = 5'h6;
assign v$C2_23_out0 = 1'h0;
assign v$C8_13_out0 = 5'h0;
assign v$ZERO_295_out0 = v$C1_2376_out0;
assign v$ZERO_296_out0 = v$C1_2377_out0;
assign v$R0_925_out0 = v$REG0_4539_out0;
assign v$R0_926_out0 = v$REG0_4540_out0;
assign v$PC1_987_out0 = v$REG1_374_out0;
assign v$PC1_988_out0 = v$REG1_375_out0;
assign v$R0_1056_out0 = v$REG0_4539_out0;
assign v$R0_1057_out0 = v$REG0_4540_out0;
assign v$C_1100_out0 = v$FF2_2554_out0;
assign v$C_1101_out0 = v$FF2_2555_out0;
assign v$R0S_1231_out0 = v$REG1_2682_out0;
assign v$R0S_1232_out0 = v$REG1_2683_out0;
assign v$EQ2_1471_out0 = v$FF1_2233_out0 == 1'h1;
assign v$Q_1495_out0 = v$FF1_2233_out0;
assign v$_1660_out0 = { v$FF3_4436_out0,v$FF4_3156_out0 };
assign v$_1661_out0 = { v$FF3_4437_out0,v$FF4_3157_out0 };
assign v$R3_1883_out0 = v$REG3_2962_out0;
assign v$R3_1884_out0 = v$REG3_2963_out0;
assign v$G11_2141_out0 = ! v$FF1_2042_out0;
assign v$G11_2142_out0 = ! v$FF1_2043_out0;
assign v$R2_2167_out0 = v$REG2_4872_out0;
assign v$R2_2168_out0 = v$REG2_4873_out0;
assign v$RAMOUT_2337_out0 = v$RAM3_1304_out0;
assign v$INTERRUPT1_2431_out0 = v$INTERRUPT1_3115_out0;
assign v$PRIORITY_2626_out0 = v$FF2_3299_out0;
assign v$PRIORITY_2627_out0 = v$FF2_3300_out0;
assign v$R3_2875_out0 = v$REG3_2962_out0;
assign v$R3_2876_out0 = v$REG3_2963_out0;
assign {v$A1_2902_out1,v$A1_2902_out0 } = v$REG1_374_out0 + v$C1_1742_out0 + v$C1_1176_out0;
assign {v$A1_2903_out1,v$A1_2903_out0 } = v$REG1_375_out0 + v$C1_1743_out0 + v$C1_1177_out0;
assign v$R2_3009_out0 = v$REG2_4872_out0;
assign v$R2_3010_out0 = v$REG2_4873_out0;
assign v$STOREDPC_3150_out0 = v$REG2_750_out0;
assign v$STOREDPC_3151_out0 = v$REG2_751_out0;
assign v$ZERO_3207_out0 = v$C1_3658_out0;
assign v$ZERO_3208_out0 = v$C1_3659_out0;
assign v$G5_3298_out0 = ! v$FF1_846_out0;
assign v$ZERO_3309_out0 = v$C1_4009_out0;
assign v$ZERO_3310_out0 = v$C1_4010_out0;
assign v$G3_3356_out0 = ! v$FF1_144_out0;
assign v$G3_3357_out0 = ! v$FF1_145_out0;
assign v$R2S_3521_out0 = v$REG3_2164_out0;
assign v$R2S_3522_out0 = v$REG3_2165_out0;
assign v$EQ1_3574_out0 = v$FF1_2233_out0 == 1'h0;
assign v$_3616_out0 = { v$FF1_1618_out0,v$FF2_4169_out0 };
assign v$_3617_out0 = { v$FF1_1619_out0,v$FF2_4170_out0 };
assign v$R1_3682_out0 = v$REG1_1399_out0;
assign v$R1_3683_out0 = v$REG1_1400_out0;
assign v$EQ2_4118_out0 = v$REG1_3272_out0 == 16'h0;
assign v$EQ2_4119_out0 = v$REG1_3273_out0 == 16'h0;
assign v$R1_4338_out0 = v$REG1_1399_out0;
assign v$R1_4339_out0 = v$REG1_1400_out0;
assign v$PC_4346_out0 = v$REG1_374_out0;
assign v$PC_4347_out0 = v$REG1_375_out0;
assign v$R3S_4759_out0 = v$REG4_1772_out0;
assign v$R3S_4760_out0 = v$REG4_1773_out0;
assign v$INTERRUPT2_4761_out0 = v$INTERRUPT2_976_out0;
assign v$1_4806_out0 = v$REG4_4843_out0[15:15];
assign v$1_4807_out0 = v$REG4_4844_out0[15:15];
assign v$FPOUT_4831_out0 = v$REG1_1106_out0;
assign v$R1S_4900_out0 = v$REG2_2762_out0;
assign v$R1S_4901_out0 = v$REG2_2763_out0;
assign v$CYC2_333_out0 = v$EQ2_1471_out0;
assign v$PRIORITYCODE_501_out0 = v$PRIORITY_2627_out0;
assign v$PRIORITYCODE_502_out0 = v$PRIORITY_2626_out0;
assign v$SEL2_1112_out0 = v$Q_1495_out0[0:0];
assign v$SHIFTPREVIOUS_1586_out0 = v$_1660_out0;
assign v$SHIFTPREVIOUS_1587_out0 = v$_1661_out0;
assign v$INTERRUPT_3178_out0 = v$INTERRUPT1_2431_out0;
assign v$INTERRUPT_3179_out0 = v$INTERRUPT2_4761_out0;
assign v$Q_3845_out0 = v$_3616_out0;
assign v$Q_3846_out0 = v$_3617_out0;
assign v$CYC1_3894_out0 = v$EQ1_3574_out0;
assign v$X_4262_out0 = v$A1_2902_out1;
assign v$X_4263_out0 = v$A1_2903_out1;
assign v$FPOUT_4289_out0 = v$FPOUT_4831_out0;
assign v$STOREDPC_5240_out0 = v$STOREDPC_3150_out0;
assign v$STOREDPC_5241_out0 = v$STOREDPC_3151_out0;
assign v$PRIORITYSAME_5355_out0 = v$G5_3298_out0;
assign v$INTERRUPT_93_out0 = v$INTERRUPT_3178_out0;
assign v$INTERRUPT_94_out0 = v$INTERRUPT_3179_out0;
assign v$G2_299_out0 = ! v$SEL2_1112_out0;
assign v$Q0_356_out0 = v$SEL2_1112_out0;
assign v$CYC2_1461_out0 = v$CYC2_333_out0;
assign v$EQ3_1928_out0 = v$SHIFTPREVIOUS_1586_out0 == 2'h2;
assign v$EQ3_1929_out0 = v$SHIFTPREVIOUS_1587_out0 == 2'h2;
assign v$EQ2_2556_out0 = v$SHIFTPREVIOUS_1586_out0 == 2'h1;
assign v$EQ2_2557_out0 = v$SHIFTPREVIOUS_1587_out0 == 2'h1;
assign v$CYC1_3443_out0 = v$CYC1_3894_out0;
assign v$EQ3_4403_out0 = v$Q_3845_out0 == 2'h2;
assign v$EQ3_4404_out0 = v$Q_3846_out0 == 2'h2;
assign v$EQ1_4689_out0 = v$Q_3845_out0 == 2'h1;
assign v$EQ1_4690_out0 = v$Q_3846_out0 == 2'h1;
assign v$EQ2_5128_out0 = v$Q_3845_out0 == 2'h0;
assign v$EQ2_5129_out0 = v$Q_3846_out0 == 2'h0;
assign v$Q_5292_out0 = v$Q_3845_out0;
assign v$Q_5293_out0 = v$Q_3846_out0;
assign v$MUX3_5300_out0 = v$FF4_89_out0 ? v$FPOUT_4289_out0 : v$RAMOUT_2337_out0;
assign v$NQ0_5_out0 = v$G2_299_out0;
assign v$DATA_968_out0 = v$MUX3_5300_out0;
assign v$_1749_out0 = v$Q_5292_out0[1:1];
assign v$_1750_out0 = v$Q_5293_out0[1:1];
assign v$G1_1924_out0 = v$EQ2_2556_out0 && v$FF2_4405_out0;
assign v$G1_1925_out0 = v$EQ2_2557_out0 && v$FF2_4406_out0;
assign v$CYC2_2652_out0 = v$CYC2_1461_out0;
assign v$FETCH_2877_out0 = v$EQ2_5128_out0;
assign v$FETCH_2878_out0 = v$EQ2_5129_out0;
assign v$EXEC1_3460_out0 = v$EQ1_4689_out0;
assign v$EXEC1_3461_out0 = v$EQ1_4690_out0;
assign v$_4077_out0 = v$Q_5292_out0[0:0];
assign v$_4078_out0 = v$Q_5293_out0[0:0];
assign v$G2_4167_out0 = v$FF1_1575_out0 && v$EQ3_1928_out0;
assign v$G2_4168_out0 = v$FF1_1576_out0 && v$EQ3_1929_out0;
assign v$EXEC2_5106_out0 = v$EQ3_4403_out0;
assign v$EXEC2_5107_out0 = v$EQ3_4404_out0;
assign v$EXEC1_201_out0 = v$EXEC1_3460_out0;
assign v$EXEC1_202_out0 = v$EXEC1_3461_out0;
assign v$CYC2_674_out0 = v$CYC2_2652_out0;
assign v$G1_909_out0 = ! v$_1749_out0;
assign v$G1_910_out0 = ! v$_1750_out0;
assign v$EXEC2_1703_out0 = v$EXEC2_5106_out0;
assign v$EXEC2_1704_out0 = v$EXEC2_5107_out0;
assign v$FETCH_2291_out0 = v$FETCH_2877_out0;
assign v$FETCH_2292_out0 = v$FETCH_2878_out0;
assign v$DMDATA_5169_out0 = v$DATA_968_out0;
assign v$EXEC2_562_out0 = v$EXEC2_1703_out0;
assign v$EXEC2_563_out0 = v$EXEC2_1704_out0;
assign v$FETCH_3722_out0 = v$FETCH_2291_out0;
assign v$FETCH_3723_out0 = v$FETCH_2292_out0;
assign v$EXEC1_3981_out0 = v$EXEC1_201_out0;
assign v$EXEC1_3982_out0 = v$EXEC1_202_out0;
assign v$DMDATA_4516_out0 = v$DMDATA_5169_out0;
assign v$FETCH_921_out0 = v$FETCH_3722_out0;
assign v$FETCH_922_out0 = v$FETCH_3723_out0;
assign v$G3_2338_out0 = v$EXEC2_562_out0 && v$FF1_4133_out0;
assign v$G3_2339_out0 = v$EXEC2_563_out0 && v$FF1_4134_out0;
assign v$EXEC1_2363_out0 = v$EXEC1_3981_out0;
assign v$EXEC1_2364_out0 = v$EXEC1_3982_out0;
assign v$READDATA1_3559_out0 = v$DMDATA_4516_out0;
assign v$READDATA2_3664_out0 = v$DMDATA_4516_out0;
assign v$EXEC2_3776_out0 = v$EXEC2_562_out0;
assign v$EXEC2_3777_out0 = v$EXEC2_563_out0;
assign v$EXEC2_4061_out0 = v$EXEC2_562_out0;
assign v$EXEC2_4062_out0 = v$EXEC2_563_out0;
assign v$EXEC1_4080_out0 = v$EXEC1_3981_out0;
assign v$EXEC1_4081_out0 = v$EXEC1_3982_out0;
assign v$G8_4101_out0 = v$EXEC2_562_out0 && v$INTERRUPT_93_out0;
assign v$G8_4102_out0 = v$EXEC2_563_out0 && v$INTERRUPT_94_out0;
assign v$G6_4510_out0 = v$INTERRUPT_93_out0 && v$FETCH_3722_out0;
assign v$G6_4511_out0 = v$INTERRUPT_94_out0 && v$FETCH_3723_out0;
assign v$G4_4743_out0 = v$INTERRUPT_93_out0 || v$FETCH_3722_out0;
assign v$G4_4744_out0 = v$INTERRUPT_94_out0 || v$FETCH_3723_out0;
assign v$G2_5045_out0 = v$FF1_4133_out0 && v$FETCH_3722_out0;
assign v$G2_5046_out0 = v$FF1_4134_out0 && v$FETCH_3723_out0;
assign v$F2_288_out0 = v$FETCH_922_out0;
assign v$EXEC2_1668_out0 = v$EXEC2_4061_out0;
assign v$EXEC2_1669_out0 = v$EXEC2_4062_out0;
assign v$READDATA1_2193_out0 = v$READDATA1_3559_out0;
assign v$EXEC2_2224_out0 = v$EXEC2_3776_out0;
assign v$EXEC2_2225_out0 = v$EXEC2_3777_out0;
assign v$G2_2236_out0 = v$EXEC1_2363_out0 && v$G3_3356_out0;
assign v$G2_2237_out0 = v$EXEC1_2364_out0 && v$G3_3357_out0;
assign v$READDATA2_2400_out0 = v$READDATA2_3664_out0;
assign v$EXEC1_3733_out0 = v$EXEC1_4080_out0;
assign v$EXEC1_3734_out0 = v$EXEC1_4081_out0;
assign v$G7_5039_out0 = v$G8_4101_out0 || v$G3_2338_out0;
assign v$G7_5040_out0 = v$G8_4102_out0 || v$G3_2339_out0;
assign v$G5_5319_out0 = v$G2_5045_out0 || v$G6_4510_out0;
assign v$G5_5320_out0 = v$G2_5046_out0 || v$G6_4511_out0;
assign v$F1_5396_out0 = v$FETCH_921_out0;
assign v$EXEC2_543_out0 = v$EXEC2_1668_out0;
assign v$EXEC2_544_out0 = v$EXEC2_1669_out0;
assign v$MUX4_936_out0 = v$FF5_271_out0 ? v$READDATA2_2400_out0 : v$ROM4_4954_out0;
assign v$MUX1_1219_out0 = v$FF2_1859_out0 ? v$READDATA1_2193_out0 : v$ROM3_3844_out0;
assign v$STORESHADOW_2370_out0 = v$G5_5319_out0;
assign v$STORESHADOW_2371_out0 = v$G5_5320_out0;
assign v$EXEC1_2956_out0 = v$EXEC1_3733_out0;
assign v$EXEC1_2957_out0 = v$EXEC1_3734_out0;
assign v$interruptatexec2_3984_out0 = v$G7_5039_out0;
assign v$interruptatexec2_3985_out0 = v$G7_5040_out0;
assign v$EXEC2_4383_out0 = v$EXEC2_1668_out0;
assign v$EXEC2_4384_out0 = v$EXEC2_1669_out0;
assign v$STORESHADOW_632_out0 = v$STORESHADOW_2370_out0;
assign v$STORESHADOW_633_out0 = v$STORESHADOW_2371_out0;
assign v$EXEC2_2321_out0 = v$EXEC2_543_out0;
assign v$EXEC2_2322_out0 = v$EXEC2_544_out0;
assign v$G10_3145_out0 = v$EXEC1_2956_out0 && v$G11_2141_out0;
assign v$G10_3146_out0 = v$EXEC1_2957_out0 && v$G11_2142_out0;
assign v$PCORROM_3465_out0 = v$MUX1_1219_out0;
assign v$PCORROM_3466_out0 = v$MUX4_936_out0;
assign v$STORESHADOW_3540_out0 = v$STORESHADOW_2370_out0;
assign v$STORESHADOW_3541_out0 = v$STORESHADOW_2371_out0;
assign v$EXEC2_4334_out0 = v$EXEC2_4383_out0;
assign v$EXEC2_4335_out0 = v$EXEC2_4384_out0;
assign v$INTERRUPT_4487_out0 = v$interruptatexec2_3984_out0;
assign v$INTERRUPT_4488_out0 = v$interruptatexec2_3985_out0;
assign v$interruptatexec2_5035_out0 = v$interruptatexec2_3984_out0;
assign v$interruptatexec2_5036_out0 = v$interruptatexec2_3985_out0;
assign v$STORESHADOW_859_out0 = v$STORESHADOW_3540_out0;
assign v$STORESHADOW_860_out0 = v$STORESHADOW_3541_out0;
assign v$STORESHADOW_1626_out0 = v$STORESHADOW_3540_out0;
assign v$STORESHADOW_1627_out0 = v$STORESHADOW_3541_out0;
assign v$STORESHADOW_1787_out0 = v$STORESHADOW_3540_out0;
assign v$STORESHADOW_1788_out0 = v$STORESHADOW_3541_out0;
assign v$RAMDOUT_2885_out0 = v$PCORROM_3465_out0;
assign v$RAMDOUT_2886_out0 = v$PCORROM_3466_out0;
assign v$STORESHADOW_3475_out0 = v$STORESHADOW_632_out0;
assign v$STORESHADOW_3476_out0 = v$STORESHADOW_633_out0;
assign v$interruptatexec2_4897_out0 = v$interruptatexec2_5035_out0;
assign v$interruptatexec2_4898_out0 = v$interruptatexec2_5036_out0;
assign v$G3_2198_out0 = v$STORESHADOW_3475_out0 || v$interruptatexec2_4897_out0;
assign v$G3_2199_out0 = v$STORESHADOW_3476_out0 || v$interruptatexec2_4898_out0;
assign v$RAMDOUT_2667_out0 = v$RAMDOUT_2885_out0;
assign v$RAMDOUT_2668_out0 = v$RAMDOUT_2886_out0;
assign v$RAMDOUT_2768_out0 = v$RAMDOUT_2885_out0;
assign v$RAMDOUT_2769_out0 = v$RAMDOUT_2886_out0;
assign v$STORESHADOW_4961_out0 = v$STORESHADOW_1787_out0;
assign v$STORESHADOW_4962_out0 = v$STORESHADOW_1788_out0;
assign v$IJUMP_1376_out0 = v$G3_2198_out0;
assign v$IJUMP_1377_out0 = v$G3_2199_out0;
assign v$MUX1_2744_out0 = v$G2_2236_out0 ? v$RAMDOUT_2667_out0 : v$REG1_3653_out0;
assign v$MUX1_2745_out0 = v$G2_2237_out0 ? v$RAMDOUT_2668_out0 : v$REG1_3654_out0;
assign v$RAMDOUT_4700_out0 = v$RAMDOUT_2768_out0;
assign v$RAMDOUT_4701_out0 = v$RAMDOUT_2769_out0;
assign v$CONTEXTSAVEN_5332_out0 = v$STORESHADOW_4961_out0;
assign v$CONTEXTSAVEN_5333_out0 = v$STORESHADOW_4962_out0;
assign v$IR_269_out0 = v$MUX1_2744_out0;
assign v$IR_270_out0 = v$MUX1_2745_out0;
assign v$RAMDOUT_2103_out0 = v$RAMDOUT_4700_out0;
assign v$RAMDOUT_2104_out0 = v$RAMDOUT_4701_out0;
assign v$_4504_out0 = v$MUX1_2744_out0[11:0];
assign v$_4504_out1 = v$MUX1_2744_out0[15:4];
assign v$_4505_out0 = v$MUX1_2745_out0[11:0];
assign v$_4505_out1 = v$MUX1_2745_out0[15:4];
assign v$EQ7_425_out0 = v$_4504_out1 == 4'h6;
assign v$EQ7_426_out0 = v$_4505_out1 == 4'h6;
assign v$EQ5_1611_out0 = v$_4504_out1 == 4'h4;
assign v$EQ5_1612_out0 = v$_4505_out1 == 4'h4;
assign v$EQ6_3613_out0 = v$_4504_out1 == 4'h5;
assign v$EQ6_3614_out0 = v$_4505_out1 == 4'h5;
assign v$EQ8_3736_out0 = v$_4504_out1 == 4'h7;
assign v$EQ8_3737_out0 = v$_4505_out1 == 4'h7;
assign v$IR110_4921_out0 = v$_4504_out0;
assign v$IR110_4922_out0 = v$_4505_out0;
assign v$IR16_5206_out0 = v$IR_269_out0;
assign v$IR16_5207_out0 = v$IR_270_out0;
assign v$EQ1_5269_out0 = v$_4504_out1 == 4'h3;
assign v$EQ1_5270_out0 = v$_4505_out1 == 4'h3;
assign v$SEL1_565_out0 = v$IR16_5206_out0[15:12];
assign v$SEL1_566_out0 = v$IR16_5207_out0[15:12];
assign v$G1_1184_out0 = v$INTERRUPT_4487_out0 || v$EQ5_1611_out0;
assign v$G1_1185_out0 = v$INTERRUPT_4488_out0 || v$EQ5_1612_out0;
assign v$SEL2_1234_out0 = v$IR16_5206_out0[9:9];
assign v$SEL2_1235_out0 = v$IR16_5207_out0[9:9];
assign v$JEQN_2145_out0 = v$EQ7_425_out0;
assign v$JEQN_2146_out0 = v$EQ7_426_out0;
assign v$STP_2446_out0 = v$EQ8_3736_out0;
assign v$STP_2447_out0 = v$EQ8_3737_out0;
assign v$JMIN_2697_out0 = v$EQ6_3613_out0;
assign v$JMIN_2698_out0 = v$EQ6_3614_out0;
assign v$IR12_3283_out0 = v$IR110_4921_out0;
assign v$IR12_3284_out0 = v$IR110_4922_out0;
assign v$IR_3909_out0 = v$IR16_5206_out0;
assign v$IR_3910_out0 = v$IR16_5207_out0;
assign v$RET_4161_out0 = v$EQ1_5269_out0;
assign v$RET_4162_out0 = v$EQ1_5270_out0;
assign v$3_31_out0 = v$IR_3909_out0[1:0];
assign v$3_32_out0 = v$IR_3910_out0[1:0];
assign v$8_112_out0 = v$IR_3909_out0[11:10];
assign v$8_113_out0 = v$IR_3910_out0[11:10];
assign v$JMIN_234_out0 = v$JMIN_2697_out0;
assign v$JMIN_235_out0 = v$JMIN_2698_out0;
assign v$JMPN_1855_out0 = v$G1_1184_out0;
assign v$JMPN_1856_out0 = v$G1_1185_out0;
assign v$IR_2357_out0 = v$IR_3909_out0;
assign v$IR_2358_out0 = v$IR_3910_out0;
assign v$EQ1_2628_out0 = v$SEL1_565_out0 == 4'h0;
assign v$EQ1_2629_out0 = v$SEL1_566_out0 == 4'h0;
assign v$JEQN_3047_out0 = v$JEQN_2145_out0;
assign v$JEQN_3048_out0 = v$JEQN_2146_out0;
assign v$7_4107_out0 = v$IR_3909_out0[15:15];
assign v$7_4108_out0 = v$IR_3910_out0[15:15];
assign v$G9_4109_out0 = v$SEL2_1234_out0 && v$EXEC1_3981_out0;
assign v$G9_4110_out0 = v$SEL2_1235_out0 && v$EXEC1_3982_out0;
assign v$RET_4312_out0 = v$RET_4161_out0;
assign v$RET_4313_out0 = v$RET_4162_out0;
assign v$1_4387_out0 = v$IR_3909_out0[14:12];
assign v$1_4388_out0 = v$IR_3910_out0[14:12];
assign v$STP_4410_out0 = v$STP_2446_out0;
assign v$STP_4411_out0 = v$STP_2447_out0;
assign v$N_5020_out0 = v$IR12_3283_out0;
assign v$N_5021_out0 = v$IR12_3284_out0;
assign v$IR15_322_out0 = v$7_4107_out0;
assign v$IR15_323_out0 = v$7_4108_out0;
assign v$5_609_out0 = v$IR_2357_out0[7:4];
assign v$5_610_out0 = v$IR_2358_out0[7:4];
assign v$RET_622_out0 = v$RET_4312_out0;
assign v$RET_623_out0 = v$RET_4313_out0;
assign v$OP_966_out0 = v$1_4387_out0;
assign v$OP_967_out0 = v$1_4388_out0;
assign v$JMPN_1036_out0 = v$JMPN_1855_out0;
assign v$JMPN_1037_out0 = v$JMPN_1856_out0;
assign v$9_1087_out0 = v$IR_2357_out0[3:2];
assign v$9_1088_out0 = v$IR_2358_out0[3:2];
assign v$M_1134_out0 = v$3_31_out0;
assign v$M_1135_out0 = v$3_32_out0;
assign v$STP_1717_out0 = v$STP_4410_out0;
assign v$STP_1718_out0 = v$STP_4411_out0;
assign v$2_1783_out0 = v$IR_2357_out0[8:8];
assign v$2_1784_out0 = v$IR_2358_out0[8:8];
assign v$G14_1860_out0 = v$INTERRUPT_93_out0 || v$RET_4312_out0;
assign v$G14_1861_out0 = v$INTERRUPT_94_out0 || v$RET_4313_out0;
assign v$RET_2021_out0 = v$RET_4312_out0;
assign v$RET_2022_out0 = v$RET_4313_out0;
assign v$4_2262_out0 = v$IR_2357_out0[4:0];
assign v$4_2263_out0 = v$IR_2358_out0[4:0];
assign v$IR_2617_out0 = v$IR_2357_out0;
assign v$IR_2618_out0 = v$IR_2358_out0;
assign v$D_2851_out0 = v$8_112_out0;
assign v$D_2852_out0 = v$8_113_out0;
assign v$MUX6_3430_out0 = v$interruptatexec2_4897_out0 ? v$C4_3093_out0 : v$N_5020_out0;
assign v$MUX6_3431_out0 = v$interruptatexec2_4898_out0 ? v$C4_3094_out0 : v$N_5021_out0;
assign v$6_4279_out0 = v$IR_2357_out0[9:9];
assign v$6_4280_out0 = v$IR_2358_out0[9:9];
assign v$G10_5141_out0 = v$EQ1_2628_out0 && v$G9_4109_out0;
assign v$G10_5142_out0 = v$EQ1_2629_out0 && v$G9_4110_out0;
assign v$K_135_out0 = v$4_2262_out0;
assign v$K_136_out0 = v$4_2263_out0;
assign v$OP_534_out0 = v$OP_966_out0;
assign v$OP_535_out0 = v$OP_967_out0;
assign v$RET_677_out0 = v$RET_622_out0;
assign v$RET_678_out0 = v$RET_623_out0;
assign v$IR_837_out0 = v$IR_2617_out0;
assign v$IR_838_out0 = v$IR_2618_out0;
assign v$C_903_out0 = v$6_4279_out0;
assign v$C_904_out0 = v$6_4280_out0;
assign v$MUX2_981_out0 = v$EXEC2_1668_out0 ? v$D_2851_out0 : v$M_1134_out0;
assign v$MUX2_982_out0 = v$EXEC2_1669_out0 ? v$D_2852_out0 : v$M_1135_out0;
assign v$JMP_2029_out0 = v$JMPN_1036_out0;
assign v$JMP_2030_out0 = v$JMPN_1037_out0;
assign v$SHIFT_2188_out0 = v$9_1087_out0;
assign v$SHIFT_2189_out0 = v$9_1088_out0;
assign v$RET_2207_out0 = v$RET_2021_out0;
assign v$RET_2208_out0 = v$RET_2022_out0;
assign v$RET_2238_out0 = v$RET_622_out0;
assign v$RET_2239_out0 = v$RET_623_out0;
assign v$IR15_2859_out0 = v$IR15_322_out0;
assign v$IR15_2860_out0 = v$IR15_323_out0;
assign v$READREQ_2930_out0 = v$G10_5141_out0;
assign v$READREQ_2931_out0 = v$G10_5142_out0;
assign v$RET_3361_out0 = v$RET_622_out0;
assign v$RET_3362_out0 = v$RET_623_out0;
assign v$B_3493_out0 = v$5_609_out0;
assign v$B_3494_out0 = v$5_610_out0;
assign v$AD2_4281_out0 = v$M_1134_out0;
assign v$AD2_4282_out0 = v$M_1135_out0;
assign v$S_4391_out0 = v$2_1783_out0;
assign v$S_4392_out0 = v$2_1784_out0;
assign v$AD1_5401_out0 = v$D_2851_out0;
assign v$AD1_5402_out0 = v$D_2852_out0;
assign v$AND_46_out0 = v$OP_534_out0 == 3'h6;
assign v$AND_47_out0 = v$OP_535_out0 == 3'h6;
assign v$G1_554_out0 = v$EXEC2_4334_out0 && v$IR15_2859_out0;
assign v$G1_555_out0 = v$EXEC2_4335_out0 && v$IR15_2860_out0;
assign v$B_578_out0 = v$B_3493_out0;
assign v$B_579_out0 = v$B_3494_out0;
assign v$TST_826_out0 = v$OP_534_out0 == 3'h7;
assign v$TST_827_out0 = v$OP_535_out0 == 3'h7;
assign v$_948_out0 = { v$K_135_out0,v$C1_1146_out0 };
assign v$_949_out0 = { v$K_136_out0,v$C1_1147_out0 };
assign v$G1_983_out0 = v$JMP_2029_out0 || v$RET_2021_out0;
assign v$G1_984_out0 = v$JMP_2030_out0 || v$RET_2022_out0;
assign v$6_998_out0 = v$IR_837_out0[1:0];
assign v$6_999_out0 = v$IR_838_out0[1:0];
assign v$C_1132_out0 = v$C_903_out0;
assign v$C_1133_out0 = v$C_904_out0;
assign v$8_1388_out0 = v$IR_837_out0[8:8];
assign v$8_1389_out0 = v$IR_838_out0[8:8];
assign v$_1879_out0 = v$AD2_4281_out0[0:0];
assign v$_1879_out1 = v$AD2_4281_out0[1:1];
assign v$_1880_out0 = v$AD2_4282_out0[0:0];
assign v$_1880_out1 = v$AD2_4282_out0[1:1];
assign v$RET_2085_out0 = v$RET_677_out0;
assign v$RET_2086_out0 = v$RET_678_out0;
assign v$7_2174_out0 = v$IR_837_out0[6:6];
assign v$7_2175_out0 = v$IR_838_out0[6:6];
assign v$4_2287_out0 = v$IR_837_out0[15:12];
assign v$4_2288_out0 = v$IR_838_out0[15:12];
assign v$3_2559_out0 = v$IR_837_out0[7:7];
assign v$3_2560_out0 = v$IR_838_out0[7:7];
assign v$9_3069_out0 = v$IR_837_out0[5:2];
assign v$9_3070_out0 = v$IR_838_out0[5:2];
assign v$ADC_3104_out0 = v$OP_534_out0 == 3'h2;
assign v$ADC_3105_out0 = v$OP_535_out0 == 3'h2;
assign v$CMP_3183_out0 = v$OP_534_out0 == 3'h5;
assign v$CMP_3184_out0 = v$OP_535_out0 == 3'h5;
assign v$_3191_out0 = v$AD1_5401_out0[0:0];
assign v$_3191_out1 = v$AD1_5401_out0[1:1];
assign v$_3192_out0 = v$AD1_5402_out0[0:0];
assign v$_3192_out1 = v$AD1_5402_out0[1:1];
assign v$S_3348_out0 = v$S_4391_out0;
assign v$S_3349_out0 = v$S_4392_out0;
assign v$SUB_3369_out0 = v$OP_534_out0 == 3'h1;
assign v$SUB_3370_out0 = v$OP_535_out0 == 3'h1;
assign v$ADD_3399_out0 = v$OP_534_out0 == 3'h0;
assign v$ADD_3400_out0 = v$OP_535_out0 == 3'h0;
assign v$2_3526_out0 = v$IR_837_out0[11:10];
assign v$2_3527_out0 = v$IR_838_out0[11:10];
assign v$MOV_3738_out0 = v$OP_534_out0 == 3'h4;
assign v$MOV_3739_out0 = v$OP_535_out0 == 3'h4;
assign v$AD3_4063_out0 = v$MUX2_981_out0;
assign v$AD3_4064_out0 = v$MUX2_982_out0;
assign v$5_4083_out0 = v$IR_837_out0[9:9];
assign v$5_4084_out0 = v$IR_838_out0[9:9];
assign v$SBC_4704_out0 = v$OP_534_out0 == 3'h3;
assign v$SBC_4705_out0 = v$OP_535_out0 == 3'h3;
assign v$SR_4826_out0 = v$SHIFT_2188_out0;
assign v$SR_4827_out0 = v$SHIFT_2189_out0;
assign v$READREQ_5066_out0 = v$READREQ_2930_out0;
assign v$READREQ_5067_out0 = v$READREQ_2931_out0;
assign v$U_54_out0 = v$7_2174_out0;
assign v$U_55_out0 = v$7_2175_out0;
assign v$G11_110_out0 = v$S_3348_out0 && v$EXEC2_4334_out0;
assign v$G11_111_out0 = v$S_3349_out0 && v$EXEC2_4335_out0;
assign v$MUX4_413_out0 = v$_1879_out0 ? v$R1_3682_out0 : v$R0_925_out0;
assign v$MUX4_414_out0 = v$_1880_out0 ? v$R1_3683_out0 : v$R0_926_out0;
assign v$D_539_out0 = v$2_3526_out0;
assign v$D_540_out0 = v$2_3527_out0;
assign v$P_905_out0 = v$3_2559_out0;
assign v$P_906_out0 = v$3_2560_out0;
assign v$B_985_out0 = v$B_578_out0;
assign v$B_986_out0 = v$B_579_out0;
assign v$CMP_1059_out0 = v$CMP_3183_out0;
assign v$CMP_1060_out0 = v$CMP_3184_out0;
assign v$TST_1125_out0 = v$TST_826_out0;
assign v$TST_1126_out0 = v$TST_827_out0;
assign v$ADC_1287_out0 = v$ADC_3104_out0;
assign v$ADC_1288_out0 = v$ADC_3105_out0;
assign v$L_1597_out0 = v$5_4083_out0;
assign v$L_1598_out0 = v$5_4084_out0;
assign v$MUX8_1725_out0 = v$RET_2085_out0 ? v$R1S_4900_out0 : v$R1_3682_out0;
assign v$MUX8_1726_out0 = v$RET_2086_out0 ? v$R1S_4901_out0 : v$R1_3683_out0;
assign v$G2_1760_out0 = v$G1_983_out0 || v$G3_2198_out0;
assign v$G2_1761_out0 = v$G1_984_out0 || v$G3_2199_out0;
assign v$W_1874_out0 = v$8_1388_out0;
assign v$W_1875_out0 = v$8_1389_out0;
assign v$MOV_1952_out0 = v$MOV_3738_out0;
assign v$MOV_1953_out0 = v$MOV_3739_out0;
assign v$SBC_2040_out0 = v$SBC_4704_out0;
assign v$SBC_2041_out0 = v$SBC_4705_out0;
assign v$MUX10_2171_out0 = v$RET_2085_out0 ? v$R3S_4759_out0 : v$R3_2875_out0;
assign v$MUX10_2172_out0 = v$RET_2086_out0 ? v$R3S_4760_out0 : v$R3_2876_out0;
assign v$AND_2179_out0 = v$AND_46_out0;
assign v$AND_2180_out0 = v$AND_47_out0;
assign v$O_2429_out0 = v$4_2287_out0;
assign v$O_2430_out0 = v$4_2288_out0;
assign v$SUB_2466_out0 = v$SUB_3369_out0;
assign v$SUB_2467_out0 = v$SUB_3370_out0;
assign v$C_2643_out0 = v$C_1132_out0;
assign v$C_2644_out0 = v$C_1133_out0;
assign v$N_2709_out0 = v$9_3069_out0;
assign v$N_2710_out0 = v$9_3070_out0;
assign v$MUX7_3001_out0 = v$RET_2085_out0 ? v$R0S_1231_out0 : v$R0_925_out0;
assign v$MUX7_3002_out0 = v$RET_2086_out0 ? v$R0S_1232_out0 : v$R0_926_out0;
assign v$RREQUEST_3720_out0 = v$READREQ_5067_out0;
assign v$RREQUEST_3721_out0 = v$READREQ_5066_out0;
assign v$MUX5_3743_out0 = v$_1879_out0 ? v$R3_2875_out0 : v$R2_2167_out0;
assign v$MUX5_3744_out0 = v$_1880_out0 ? v$R3_2876_out0 : v$R2_2168_out0;
assign v$MUX9_3795_out0 = v$RET_2085_out0 ? v$R2S_3521_out0 : v$R2_2167_out0;
assign v$MUX9_3796_out0 = v$RET_2086_out0 ? v$R2S_3522_out0 : v$R2_2168_out0;
assign v$M_4607_out0 = v$6_998_out0;
assign v$M_4608_out0 = v$6_999_out0;
assign v$ADD_4927_out0 = v$ADD_3399_out0;
assign v$ADD_4928_out0 = v$ADD_3400_out0;
assign v$_5317_out0 = v$B_578_out0[0:0];
assign v$_5317_out1 = v$B_578_out0[3:3];
assign v$_5318_out0 = v$B_579_out0[0:0];
assign v$_5318_out1 = v$B_579_out0[3:3];
assign v$MUX1_17_out0 = v$C_2643_out0 ? v$ROR_3251_out0 : v$SR_4826_out0;
assign v$MUX1_18_out0 = v$C_2644_out0 ? v$ROR_3252_out0 : v$SR_4827_out0;
assign v$R1S_279_out0 = v$MUX8_1725_out0;
assign v$R1S_280_out0 = v$MUX8_1726_out0;
assign v$G6_410_out0 = v$EXEC1_2956_out0 && v$W_1874_out0;
assign v$G6_411_out0 = v$EXEC1_2957_out0 && v$W_1875_out0;
assign v$EQ1_737_out0 = v$O_2429_out0 == 4'h6;
assign v$EQ1_738_out0 = v$O_2430_out0 == 4'h6;
assign v$G8_1121_out0 = v$SUB_2466_out0 || v$CMP_1059_out0;
assign v$G8_1122_out0 = v$SUB_2467_out0 || v$CMP_1060_out0;
assign v$R0S_1142_out0 = v$MUX7_3001_out0;
assign v$R0S_1143_out0 = v$MUX7_3002_out0;
assign v$R2S_1379_out0 = v$MUX9_3795_out0;
assign v$R2S_1380_out0 = v$MUX9_3796_out0;
assign v$MUX6_1469_out0 = v$_1879_out1 ? v$MUX5_3743_out0 : v$MUX4_413_out0;
assign v$MUX6_1470_out0 = v$_1880_out1 ? v$MUX5_3744_out0 : v$MUX4_414_out0;
assign v$MUX2_1594_out0 = v$ADD_4927_out0 ? v$C2_3074_out0 : v$FF1_2975_out0;
assign v$MUX2_1595_out0 = v$ADD_4928_out0 ? v$C2_3075_out0 : v$FF1_2976_out0;
assign v$U_1679_out0 = v$U_54_out0;
assign v$U_1680_out0 = v$U_55_out0;
assign v$G5_1876_out0 = ! v$MOV_1952_out0;
assign v$G5_1877_out0 = ! v$MOV_1953_out0;
assign v$B_1966_out0 = v$B_985_out0;
assign v$B_1967_out0 = v$B_986_out0;
assign v$R3TEST_2015_out0 = v$MUX10_2171_out0;
assign v$R3TEST_2016_out0 = v$MUX10_2172_out0;
assign v$_2747_out0 = v$_5317_out1[0:0];
assign v$_2747_out1 = v$_5317_out1[2:2];
assign v$_2748_out0 = v$_5318_out1[0:0];
assign v$_2748_out1 = v$_5318_out1[2:2];
assign v$EQ4_2879_out0 = v$O_2429_out0 == 4'h0;
assign v$EQ4_2880_out0 = v$O_2430_out0 == 4'h0;
assign v$G2_2927_out0 = ! v$C_2643_out0;
assign v$G2_2928_out0 = ! v$C_2644_out0;
assign v$G3_3253_out0 = v$EXEC2_2321_out0 && v$L_1597_out0;
assign v$G3_3254_out0 = v$EXEC2_2322_out0 && v$L_1598_out0;
assign v$G2_3352_out0 = ! v$L_1597_out0;
assign v$G2_3353_out0 = ! v$L_1598_out0;
assign v$EQ1_3645_out0 = v$B_985_out0 == 4'h0;
assign v$EQ1_3646_out0 = v$B_986_out0 == 4'h0;
assign v$G9_3695_out0 = !(v$CMP_1059_out0 || v$TST_1125_out0);
assign v$G9_3696_out0 = !(v$CMP_1060_out0 || v$TST_1126_out0);
assign v$G2_3757_out0 = v$SUB_2466_out0 || v$SBC_2040_out0;
assign v$G2_3758_out0 = v$SUB_2467_out0 || v$SBC_2041_out0;
assign v$EQ3_4099_out0 = v$O_2429_out0 == 4'h5;
assign v$EQ3_4100_out0 = v$O_2430_out0 == 4'h5;
assign v$G3_4378_out0 = v$ADD_4927_out0 || v$ADC_1287_out0;
assign v$G3_4379_out0 = v$ADD_4928_out0 || v$ADC_1288_out0;
assign v$R3S_4764_out0 = v$MUX10_2171_out0;
assign v$R3S_4765_out0 = v$MUX10_2172_out0;
assign v$G8_4860_out0 = v$L_1597_out0 && v$EXEC2_2321_out0;
assign v$G8_4861_out0 = v$L_1598_out0 && v$EXEC2_2322_out0;
assign v$N_5197_out0 = v$N_2709_out0;
assign v$N_5198_out0 = v$N_2710_out0;
assign v$G12_5243_out0 = v$AND_2179_out0 || v$TST_1125_out0;
assign v$G12_5244_out0 = v$AND_2180_out0 || v$TST_1126_out0;
assign v$DOUT2_1013_out0 = v$MUX6_1469_out0;
assign v$DOUT2_1014_out0 = v$MUX6_1470_out0;
assign v$EQ1_1314_out0 = v$B_1966_out0 == 4'h0;
assign v$EQ1_1315_out0 = v$B_1967_out0 == 4'h0;
assign v$EN_1424_out0 = v$_2747_out0;
assign v$EN_1425_out0 = v$_2748_out0;
assign v$MUX1_1624_out0 = v$_3191_out0 ? v$R1S_279_out0 : v$R0S_1142_out0;
assign v$MUX1_1625_out0 = v$_3192_out0 ? v$R1S_280_out0 : v$R0S_1143_out0;
assign v$G1_1886_out0 = v$EQ1_737_out0 && v$EQ2_4118_out0;
assign v$G1_1887_out0 = v$EQ1_738_out0 && v$EQ2_4119_out0;
assign v$R0TEST_2264_out0 = v$R0S_1142_out0;
assign v$R0TEST_2265_out0 = v$R0S_1143_out0;
assign v$_2484_out0 = { v$N_5197_out0,v$C1_2031_out0 };
assign v$_2485_out0 = { v$N_5198_out0,v$C1_2032_out0 };
assign v$MUX2_2857_out0 = v$_3191_out0 ? v$R3S_4764_out0 : v$R2S_1379_out0;
assign v$MUX2_2858_out0 = v$_3192_out0 ? v$R3S_4765_out0 : v$R2S_1380_out0;
assign v$SR_3148_out0 = v$MUX1_17_out0;
assign v$SR_3149_out0 = v$MUX1_18_out0;
assign v$NOR_3258_out0 = v$G9_3695_out0;
assign v$NOR_3259_out0 = v$G9_3696_out0;
assign v$MUX2_3319_out0 = v$U_1679_out0 ? v$C3_4001_out0 : v$C4_1217_out0;
assign v$MUX2_3320_out0 = v$U_1680_out0 ? v$C3_4002_out0 : v$C4_1218_out0;
assign v$G5_3518_out0 = v$G6_410_out0 || v$G3_3253_out0;
assign v$G5_3519_out0 = v$G6_411_out0 || v$G3_3254_out0;
assign v$G1_3741_out0 = v$G2_2927_out0 && v$_5317_out0;
assign v$G1_3742_out0 = v$G2_2928_out0 && v$_5318_out0;
assign v$R1TEST_4069_out0 = v$R1S_279_out0;
assign v$R1TEST_4070_out0 = v$R1S_280_out0;
assign v$_4236_out0 = v$_2747_out1[0:0];
assign v$_4236_out1 = v$_2747_out1[1:1];
assign v$_4237_out0 = v$_2748_out1[0:0];
assign v$_4237_out1 = v$_2748_out1[1:1];
assign v$G4_4284_out0 = v$1_4806_out0 && v$EQ3_4099_out0;
assign v$G4_4285_out0 = v$1_4807_out0 && v$EQ3_4100_out0;
assign v$R2TEST_4286_out0 = v$R2S_1379_out0;
assign v$R2TEST_4287_out0 = v$R2S_1380_out0;
assign v$MUX3_4659_out0 = v$G8_1121_out0 ? v$C1_3797_out0 : v$MUX2_1594_out0;
assign v$MUX3_4660_out0 = v$G8_1122_out0 ? v$C1_3798_out0 : v$MUX2_1595_out0;
assign v$G7_4776_out0 = v$G2_3757_out0 || v$CMP_1059_out0;
assign v$G7_4777_out0 = v$G2_3758_out0 || v$CMP_1060_out0;
assign v$G9_5174_out0 = v$EXEC2_2321_out0 && v$G2_3352_out0;
assign v$G9_5175_out0 = v$EXEC2_2322_out0 && v$G2_3353_out0;
assign v$R3TEST_5310_out0 = v$R3TEST_2015_out0;
assign v$R3TEST_5311_out0 = v$R3TEST_2016_out0;
assign v$WENLDST_334_out0 = v$G5_3518_out0;
assign v$WENLDST_335_out0 = v$G5_3519_out0;
assign v$MUX3_366_out0 = v$_3191_out1 ? v$MUX2_2857_out0 : v$MUX1_1624_out0;
assign v$MUX3_367_out0 = v$_3192_out1 ? v$MUX2_2858_out0 : v$MUX1_1625_out0;
assign v$SR_911_out0 = v$SR_3148_out0;
assign v$SR_912_out0 = v$SR_3149_out0;
assign v$R2TEST_1284_out0 = v$R2TEST_4286_out0;
assign v$R2TEST_1285_out0 = v$R2TEST_4287_out0;
assign v$SHIFT_1565_out0 = v$SR_3148_out0;
assign v$SHIFT_1566_out0 = v$SR_3149_out0;
assign v$XOR1_2094_out0 = v$_2484_out0 ^ v$C2_5403_out0;
assign v$XOR1_2095_out0 = v$_2485_out0 ^ v$C2_5404_out0;
assign v$G10_2259_out0 = v$G1_554_out0 && v$NOR_3258_out0;
assign v$G10_2260_out0 = v$G1_555_out0 && v$NOR_3259_out0;
assign v$SR_2469_out0 = v$SR_3148_out0;
assign v$SR_2470_out0 = v$SR_3149_out0;
assign v$R1TEST_2942_out0 = v$R1TEST_4069_out0;
assign v$R1TEST_2943_out0 = v$R1TEST_4070_out0;
assign v$CIN_3082_out0 = v$MUX3_4659_out0;
assign v$CIN_3083_out0 = v$MUX3_4660_out0;
assign v$MUX4_3084_out0 = v$RET_3361_out0 ? v$REG2_1904_out0 : v$G1_1886_out0;
assign v$MUX4_3085_out0 = v$RET_3362_out0 ? v$REG2_1905_out0 : v$G1_1887_out0;
assign v$EN_3825_out0 = v$G1_3741_out0;
assign v$EN_3826_out0 = v$G1_3742_out0;
assign v$SR_3994_out0 = v$SR_3148_out0;
assign v$SR_3995_out0 = v$SR_3149_out0;
assign v$MUX1_4052_out0 = v$G7_4776_out0 ? v$C4_395_out0 : v$C3_1545_out0;
assign v$MUX1_4053_out0 = v$G7_4777_out0 ? v$C4_396_out0 : v$C3_1546_out0;
assign v$SR_4135_out0 = v$SR_3148_out0;
assign v$SR_4136_out0 = v$SR_3149_out0;
assign v$G4_4501_out0 = v$G7_4776_out0 || v$G3_4378_out0;
assign v$G4_4502_out0 = v$G7_4777_out0 || v$G3_4379_out0;
assign v$RM_4530_out0 = v$DOUT2_1013_out0;
assign v$RM_4531_out0 = v$DOUT2_1014_out0;
assign v$MUX2_4845_out0 = v$RET_3361_out0 ? v$REG3_574_out0 : v$G4_4284_out0;
assign v$MUX2_4846_out0 = v$RET_3362_out0 ? v$REG3_575_out0 : v$G4_4285_out0;
assign v$EN_4955_out0 = v$_4236_out0;
assign v$EN_4956_out0 = v$_4237_out0;
assign v$RM_5033_out0 = v$DOUT2_1013_out0;
assign v$RM_5034_out0 = v$DOUT2_1014_out0;
assign v$R3_5058_out0 = v$R3TEST_5310_out0;
assign v$R3_5059_out0 = v$R3TEST_5311_out0;
assign v$R0TEST_5113_out0 = v$R0TEST_2264_out0;
assign v$R0TEST_5114_out0 = v$R0TEST_2265_out0;
assign v$G7_5185_out0 = v$EQ4_2879_out0 && v$G9_5174_out0;
assign v$G7_5186_out0 = v$EQ4_2880_out0 && v$G9_5175_out0;
assign v$EN_5416_out0 = v$_4236_out1;
assign v$EN_5417_out0 = v$_4237_out1;
assign v$_523_out0 = v$SR_4135_out0[0:0];
assign v$_523_out1 = v$SR_4135_out0[1:1];
assign v$_524_out0 = v$SR_4136_out0[0:0];
assign v$_524_out1 = v$SR_4136_out0[1:1];
assign v$DOUT1_873_out0 = v$MUX3_366_out0;
assign v$DOUT1_874_out0 = v$MUX3_367_out0;
assign v$EQ_923_out0 = v$MUX4_3084_out0;
assign v$EQ_924_out0 = v$MUX4_3085_out0;
assign v$WENLDST_1028_out0 = v$WENLDST_334_out0;
assign v$WENLDST_1029_out0 = v$WENLDST_335_out0;
assign v$_1244_out0 = v$SR_911_out0[0:0];
assign v$_1244_out1 = v$SR_911_out0[1:1];
assign v$_1245_out0 = v$SR_912_out0[0:0];
assign v$_1245_out1 = v$SR_912_out0[1:1];
assign v$_1569_out0 = v$SHIFT_1565_out0[0:0];
assign v$_1569_out1 = v$SHIFT_1565_out0[1:1];
assign v$_1570_out0 = v$SHIFT_1566_out0[0:0];
assign v$_1570_out1 = v$SHIFT_1566_out0[1:1];
assign v$RM_1744_out0 = v$RM_5033_out0;
assign v$RM_1745_out0 = v$RM_5034_out0;
assign v$_2186_out0 = v$SR_2469_out0[0:0];
assign v$_2186_out1 = v$SR_2469_out0[1:1];
assign v$_2187_out0 = v$SR_2470_out0[0:0];
assign v$_2187_out1 = v$SR_2470_out0[1:1];
assign v$R3_2227_out0 = v$R3_5058_out0;
assign v$R3_2228_out0 = v$R3_5059_out0;
assign v$G6_2973_out0 = v$G4_4501_out0 && v$G5_1876_out0;
assign v$G6_2974_out0 = v$G4_4502_out0 && v$G5_1877_out0;
assign v$RM_3021_out0 = v$RM_5033_out0;
assign v$RM_3022_out0 = v$RM_5034_out0;
assign v$MUX1_3023_out0 = v$U_1679_out0 ? v$_2484_out0 : v$XOR1_2094_out0;
assign v$MUX1_3024_out0 = v$U_1680_out0 ? v$_2485_out0 : v$XOR1_2095_out0;
assign v$MI_3185_out0 = v$MUX2_4845_out0;
assign v$MI_3186_out0 = v$MUX2_4846_out0;
assign v$RAMWEN_3187_out0 = v$G7_5185_out0;
assign v$RAMWEN_3188_out0 = v$G7_5186_out0;
assign v$MUX1_3674_out0 = v$C_1132_out0 ? v$_948_out0 : v$RM_4530_out0;
assign v$MUX1_3675_out0 = v$C_1133_out0 ? v$_949_out0 : v$RM_4531_out0;
assign v$_3782_out0 = v$SR_3994_out0[0:0];
assign v$_3782_out1 = v$SR_3994_out0[1:1];
assign v$_3783_out0 = v$SR_3995_out0[0:0];
assign v$_3783_out1 = v$SR_3995_out0[1:1];
assign v$R2_3953_out0 = v$R2TEST_1284_out0;
assign v$R2_3954_out0 = v$R2TEST_1285_out0;
assign v$R1_4116_out0 = v$R1TEST_2942_out0;
assign v$R1_4117_out0 = v$R1TEST_2943_out0;
assign v$R0_4215_out0 = v$R0TEST_5113_out0;
assign v$R0_4216_out0 = v$R0TEST_5114_out0;
assign v$WENALU_5353_out0 = v$G10_2259_out0;
assign v$WENALU_5354_out0 = v$G10_2260_out0;
assign v$EQ_1529_out0 = v$EQ_923_out0;
assign v$EQ_1530_out0 = v$EQ_924_out0;
assign v$R3_2053_out0 = v$R3_2227_out0;
assign v$R3_2054_out0 = v$R3_2228_out0;
assign v$RD_2135_out0 = v$DOUT1_873_out0;
assign v$RD_2136_out0 = v$DOUT1_874_out0;
assign v$RM_2274_out0 = v$RM_1744_out0;
assign v$RM_2275_out0 = v$RM_1745_out0;
assign v$SHIFTIN_2366_out0 = v$MUX1_3674_out0;
assign v$SHIFTIN_2367_out0 = v$MUX1_3675_out0;
assign v$WENALU_2753_out0 = v$WENALU_5353_out0;
assign v$WENALU_2754_out0 = v$WENALU_5354_out0;
assign v$R1_2934_out0 = v$R1_4116_out0;
assign v$R1_2935_out0 = v$R1_4117_out0;
assign v$MUX5_3080_out0 = v$G10_3145_out0 ? v$RM_3021_out0 : v$REG5_3036_out0;
assign v$MUX5_3081_out0 = v$G10_3146_out0 ? v$RM_3022_out0 : v$REG5_3037_out0;
assign v$R0_3873_out0 = v$R0_4215_out0;
assign v$R0_3874_out0 = v$R0_4216_out0;
assign v$MI_4847_out0 = v$MI_3185_out0;
assign v$MI_4848_out0 = v$MI_3186_out0;
assign v$R2_5037_out0 = v$R2_3953_out0;
assign v$R2_5038_out0 = v$R2_3954_out0;
assign v$WENRAM_5126_out0 = v$RAMWEN_3187_out0;
assign v$WENRAM_5127_out0 = v$RAMWEN_3188_out0;
assign v$RM_1148_out0 = v$MUX5_3080_out0;
assign v$RM_1149_out0 = v$MUX5_3081_out0;
assign v$MI_1295_out0 = v$MI_4847_out0;
assign v$MI_1296_out0 = v$MI_4848_out0;
assign v$RDOUT_1775_out0 = v$RD_2135_out0;
assign v$RDOUT_1776_out0 = v$RD_2136_out0;
assign v$IN_1798_out0 = v$SHIFTIN_2366_out0;
assign v$IN_1799_out0 = v$SHIFTIN_2367_out0;
assign v$WRITEREQ_2132_out0 = v$WENRAM_5126_out0;
assign v$WRITEREQ_2133_out0 = v$WENRAM_5127_out0;
assign v$R31_2229_out0 = v$R3_2053_out0;
assign v$EQ_2306_out0 = v$EQ_1529_out0;
assign v$EQ_2307_out0 = v$EQ_1530_out0;
assign v$R2_2904_out0 = v$R2_5037_out0;
assign v$R2_2905_out0 = v$R2_5038_out0;
assign v$R32_3176_out0 = v$R3_2054_out0;
assign v$R0_3907_out0 = v$R0_3873_out0;
assign v$R0_3908_out0 = v$R0_3874_out0;
assign v$OP1_4087_out0 = v$RD_2135_out0;
assign v$OP1_4088_out0 = v$RD_2136_out0;
assign v$MUX3_4875_out0 = v$IR15_322_out0 ? v$WENALU_2753_out0 : v$WENLDST_1028_out0;
assign v$MUX3_4876_out0 = v$IR15_323_out0 ? v$WENALU_2754_out0 : v$WENLDST_1029_out0;
assign v$IN_4895_out0 = v$SHIFTIN_2366_out0;
assign v$IN_4896_out0 = v$SHIFTIN_2367_out0;
assign v$R1_5052_out0 = v$R1_2934_out0;
assign v$R1_5053_out0 = v$R1_2935_out0;
assign v$RDOUT_289_out0 = v$RDOUT_1775_out0;
assign v$RDOUT_290_out0 = v$RDOUT_1776_out0;
assign v$WEN3_931_out0 = v$MUX3_4875_out0;
assign v$WEN3_932_out0 = v$MUX3_4876_out0;
assign v$OP1_1525_out0 = v$OP1_4087_out0;
assign v$OP1_1526_out0 = v$OP1_4088_out0;
assign v$MI_1823_out0 = v$MI_1295_out0;
assign v$MI_1824_out0 = v$MI_1296_out0;
assign v$R22_2273_out0 = v$R2_2905_out0;
assign v$R02_2546_out0 = v$R0_3908_out0;
assign v$R21_2715_out0 = v$R2_2904_out0;
assign v$IN_2966_out0 = v$IN_4895_out0;
assign v$IN_2967_out0 = v$IN_4896_out0;
assign v$MUX3_3233_out0 = v$EQ1_3645_out0 ? v$IN_1798_out0 : v$C1_864_out0;
assign v$MUX3_3234_out0 = v$EQ1_3646_out0 ? v$IN_1799_out0 : v$C1_865_out0;
assign v$EQ_3344_out0 = v$EQ_2306_out0;
assign v$EQ_3345_out0 = v$EQ_2307_out0;
assign v$R11_3434_out0 = v$R1_5052_out0;
assign v$RM_3453_out0 = v$RM_1148_out0;
assign v$RM_3454_out0 = v$RM_1149_out0;
assign v$R01_3542_out0 = v$R0_3907_out0;
assign v$WRITEREQ_4482_out0 = v$WRITEREQ_2132_out0;
assign v$WRITEREQ_4483_out0 = v$WRITEREQ_2133_out0;
assign v$R12_4500_out0 = v$R1_5053_out0;
assign v$WREQUEST_508_out0 = v$WRITEREQ_4483_out0;
assign v$WREQUEST_509_out0 = v$WRITEREQ_4482_out0;
assign v$_880_out0 = v$IN_2966_out0[0:0];
assign v$_880_out1 = v$IN_2966_out0[15:15];
assign v$_881_out0 = v$IN_2967_out0[0:0];
assign v$_881_out1 = v$IN_2967_out0[15:15];
assign v$WDATA_964_out0 = v$RDOUT_289_out0;
assign v$WDATA_965_out0 = v$RDOUT_290_out0;
assign {v$A1_1123_out1,v$A1_1123_out0 } = v$RM_3453_out0 + v$MUX1_3023_out0 + v$MUX2_3319_out0;
assign {v$A1_1124_out1,v$A1_1124_out0 } = v$RM_3454_out0 + v$MUX1_3024_out0 + v$MUX2_3320_out0;
assign v$G6_1567_out0 = v$EQ_3344_out0 || v$MI_1823_out0;
assign v$G6_1568_out0 = v$EQ_3345_out0 || v$MI_1824_out0;
assign v$G4_2282_out0 = v$EQ_3344_out0 || v$IJUMP_1376_out0;
assign v$G4_2283_out0 = v$EQ_3345_out0 || v$IJUMP_1377_out0;
assign v$IN_2394_out0 = v$MUX3_3233_out0;
assign v$IN_2395_out0 = v$MUX3_3234_out0;
assign v$_3534_out0 = v$IN_2966_out0[14:0];
assign v$_3534_out1 = v$IN_2966_out0[15:1];
assign v$_3535_out0 = v$IN_2967_out0[14:0];
assign v$_3535_out1 = v$IN_2967_out0[15:1];
assign v$D1_3759_out0 = (v$AD3_4063_out0 == 2'b00) ? v$WEN3_931_out0 : 1'h0;
assign v$D1_3759_out1 = (v$AD3_4063_out0 == 2'b01) ? v$WEN3_931_out0 : 1'h0;
assign v$D1_3759_out2 = (v$AD3_4063_out0 == 2'b10) ? v$WEN3_931_out0 : 1'h0;
assign v$D1_3759_out3 = (v$AD3_4063_out0 == 2'b11) ? v$WEN3_931_out0 : 1'h0;
assign v$D1_3760_out0 = (v$AD3_4064_out0 == 2'b00) ? v$WEN3_932_out0 : 1'h0;
assign v$D1_3760_out1 = (v$AD3_4064_out0 == 2'b01) ? v$WEN3_932_out0 : 1'h0;
assign v$D1_3760_out2 = (v$AD3_4064_out0 == 2'b10) ? v$WEN3_932_out0 : 1'h0;
assign v$D1_3760_out3 = (v$AD3_4064_out0 == 2'b11) ? v$WEN3_932_out0 : 1'h0;
assign v$A_4810_out0 = v$OP1_1525_out0;
assign v$A_4811_out0 = v$OP1_1526_out0;
assign v$G5_5029_out0 = v$MI_1823_out0 || v$IJUMP_1376_out0;
assign v$G5_5030_out0 = v$MI_1824_out0 || v$IJUMP_1377_out0;
assign v$_220_out0 = { v$_880_out1,v$_880_out0 };
assign v$_221_out0 = { v$_881_out1,v$_881_out0 };
assign v$WRITEDATA_1247_out0 = v$WDATA_965_out0;
assign v$WRITEDATA_1248_out0 = v$WDATA_964_out0;
assign v$MUX17_1733_out0 = v$RET_2085_out0 ? v$C1_1229_out0 : v$D1_3759_out2;
assign v$MUX17_1734_out0 = v$RET_2086_out0 ? v$C1_1230_out0 : v$D1_3760_out2;
assign v$_1816_out0 = { v$_880_out1,v$_3534_out1 };
assign v$_1817_out0 = { v$_881_out1,v$_3535_out1 };
assign v$IN_2403_out0 = v$IN_2394_out0;
assign v$IN_2404_out0 = v$IN_2395_out0;
assign v$G8_2713_out0 = v$G4_2282_out0 || v$G5_5029_out0;
assign v$G8_2714_out0 = v$G4_2283_out0 || v$G5_5030_out0;
assign v$_3045_out0 = { v$_880_out1,v$C2_620_out0 };
assign v$_3046_out0 = { v$_881_out1,v$C2_621_out0 };
assign v$RMN_3404_out0 = v$A1_1123_out0;
assign v$RMN_3405_out0 = v$A1_1124_out0;
assign v$_3799_out0 = { v$C1_5097_out0,v$_3534_out0 };
assign v$_3800_out0 = { v$C1_5098_out0,v$_3535_out0 };
assign v$G1_3963_out0 = ((v$WREQUEST_508_out0 && !v$RREQUEST_3720_out0) || (!v$WREQUEST_508_out0) && v$RREQUEST_3720_out0);
assign v$G1_3964_out0 = ((v$WREQUEST_509_out0 && !v$RREQUEST_3721_out0) || (!v$WREQUEST_509_out0) && v$RREQUEST_3721_out0);
assign v$MUX16_3996_out0 = v$RET_2085_out0 ? v$C1_1229_out0 : v$D1_3759_out1;
assign v$MUX16_3997_out0 = v$RET_2086_out0 ? v$C1_1230_out0 : v$D1_3760_out1;
assign v$MUX7_4351_out0 = v$G6_1567_out0 ? v$N_5020_out0 : v$A1_2902_out0;
assign v$MUX7_4352_out0 = v$G6_1568_out0 ? v$N_5021_out0 : v$A1_2903_out0;
assign v$MUX15_4624_out0 = v$RET_2085_out0 ? v$C1_1229_out0 : v$D1_3759_out0;
assign v$MUX15_4625_out0 = v$RET_2086_out0 ? v$C1_1230_out0 : v$D1_3760_out0;
assign v$_4906_out0 = v$A_4810_out0[0:0];
assign v$_4906_out1 = v$A_4810_out0[15:15];
assign v$_4907_out0 = v$A_4811_out0[0:0];
assign v$_4907_out1 = v$A_4811_out0[15:15];
assign v$NOTUSED_4919_out0 = v$A1_1123_out1;
assign v$NOTUSED_4920_out0 = v$A1_1124_out1;
assign v$MUX18_5025_out0 = v$RET_2085_out0 ? v$C1_1229_out0 : v$D1_3759_out3;
assign v$MUX18_5026_out0 = v$RET_2086_out0 ? v$C1_1230_out0 : v$D1_3760_out3;
assign v$_116_out0 = { v$G1_3963_out0,v$PRIORITYCODE_501_out0 };
assign v$_117_out0 = { v$G1_3964_out0,v$PRIORITYCODE_502_out0 };
assign v$ASR_628_out0 = v$_1816_out0;
assign v$ASR_629_out0 = v$_1817_out0;
assign v$RMN_844_out0 = v$RMN_3404_out0;
assign v$RMN_845_out0 = v$RMN_3405_out0;
assign v$ROR_1686_out0 = v$_220_out0;
assign v$ROR_1687_out0 = v$_221_out0;
assign v$_1728_out0 = v$_4906_out1[0:0];
assign v$_1728_out1 = v$_4906_out1[14:14];
assign v$_1729_out0 = v$_4907_out1[0:0];
assign v$_1729_out1 = v$_4907_out1[14:14];
assign v$_2284_out0 = v$IN_2403_out0[14:0];
assign v$_2284_out1 = v$IN_2403_out0[15:1];
assign v$_2285_out0 = v$IN_2404_out0[14:0];
assign v$_2285_out1 = v$IN_2404_out0[15:1];
assign v$_3772_out0 = v$IN_2403_out0[0:0];
assign v$_3772_out1 = v$IN_2403_out0[15:15];
assign v$_3773_out0 = v$IN_2404_out0[0:0];
assign v$_3773_out1 = v$IN_2404_out0[15:15];
assign v$LSL_3834_out0 = v$_3799_out0;
assign v$LSL_3835_out0 = v$_3800_out0;
assign v$G7_4011_out0 = v$G2_1760_out0 || v$G8_2713_out0;
assign v$G7_4012_out0 = v$G2_1761_out0 || v$G8_2714_out0;
assign v$LSR_4948_out0 = v$_3045_out0;
assign v$LSR_4949_out0 = v$_3046_out0;
assign v$MUX3_462_out0 = v$_3782_out1 ? v$ROR_1686_out0 : v$LSR_4948_out0;
assign v$MUX3_463_out0 = v$_3783_out1 ? v$ROR_1687_out0 : v$LSR_4949_out0;
assign v$_593_out0 = { v$G1_1924_out0,v$_2284_out0 };
assign v$_594_out0 = { v$G1_1925_out0,v$_2285_out0 };
assign v$MUX2_769_out0 = v$G7_4011_out0 ? v$MUX6_3430_out0 : v$A1_2902_out0;
assign v$MUX2_770_out0 = v$G7_4012_out0 ? v$MUX6_3431_out0 : v$A1_2903_out0;
assign v$_1238_out0 = v$_1728_out1[0:0];
assign v$_1238_out1 = v$_1728_out1[13:13];
assign v$_1239_out0 = v$_1729_out1[0:0];
assign v$_1239_out1 = v$_1729_out1[13:13];
assign v$MUX2_2109_out0 = v$_3782_out1 ? v$ASR_628_out0 : v$LSL_3834_out0;
assign v$MUX2_2110_out0 = v$_3783_out1 ? v$ASR_629_out0 : v$LSL_3835_out0;
assign v$CONTROLREQUEST_2332_out0 = v$_116_out0;
assign v$CONTROLREQUEST_2333_out0 = v$_117_out0;
assign v$MUX3_3333_out0 = v$G8_4860_out0 ? v$RAMDOUT_2103_out0 : v$RMN_844_out0;
assign v$MUX3_3334_out0 = v$G8_4861_out0 ? v$RAMDOUT_2104_out0 : v$RMN_845_out0;
assign v$MUX1_3811_out0 = v$P_905_out0 ? v$RMN_844_out0 : v$RM_1148_out0;
assign v$MUX1_3812_out0 = v$P_906_out0 ? v$RMN_845_out0 : v$RM_1149_out0;
assign v$_5287_out0 = { v$_3772_out1,v$G2_4167_out0 };
assign v$_5288_out0 = { v$_3773_out1,v$G2_4168_out0 };
assign v$MUX4_407_out0 = v$_3782_out0 ? v$MUX3_462_out0 : v$MUX2_2109_out0;
assign v$MUX4_408_out0 = v$_3783_out0 ? v$MUX3_463_out0 : v$MUX2_2110_out0;
assign v$MSL_591_out0 = v$_593_out0;
assign v$MSL_592_out0 = v$_594_out0;
assign v$MUX4_788_out0 = v$STP_1717_out0 ? v$PC_4346_out0 : v$MUX2_769_out0;
assign v$MUX4_789_out0 = v$STP_1718_out0 ? v$PC_4347_out0 : v$MUX2_770_out0;
assign v$CONTROLREQUEST1_1141_out0 = v$CONTROLREQUEST_2333_out0;
assign v$MSR_2502_out0 = v$_5287_out0;
assign v$MSR_2503_out0 = v$_5288_out0;
assign v$EA_2692_out0 = v$MUX1_3811_out0;
assign v$EA_2693_out0 = v$MUX1_3812_out0;
assign v$_3126_out0 = v$_1238_out1[0:0];
assign v$_3126_out1 = v$_1238_out1[12:12];
assign v$_3127_out0 = v$_1239_out1[0:0];
assign v$_3127_out1 = v$_1239_out1[12:12];
assign v$_3346_out0 = v$MUX1_3811_out0[11:0];
assign v$_3346_out1 = v$MUX1_3811_out0[15:4];
assign v$_3347_out0 = v$MUX1_3812_out0[11:0];
assign v$_3347_out1 = v$MUX1_3812_out0[15:4];
assign v$REGDIN_3350_out0 = v$MUX3_3333_out0;
assign v$REGDIN_3351_out0 = v$MUX3_3334_out0;
assign v$CONTROLREQUEST2_4145_out0 = v$CONTROLREQUEST_2332_out0;
assign v$ControlRequest1_214_out0 = v$CONTROLREQUEST1_1141_out0;
assign v$MUX4_276_out0 = v$_1569_out0 ? v$IN_2403_out0 : v$MSR_2502_out0;
assign v$MUX4_277_out0 = v$_1570_out0 ? v$IN_2404_out0 : v$MSR_2503_out0;
assign v$MUX1_1435_out0 = v$EN_3825_out0 ? v$MUX4_407_out0 : v$IN_2966_out0;
assign v$MUX1_1436_out0 = v$EN_3826_out0 ? v$MUX4_408_out0 : v$IN_2967_out0;
assign v$RAMADDRMUX_1479_out0 = v$_3346_out0;
assign v$RAMADDRMUX_1480_out0 = v$_3347_out0;
assign v$REGDIN_1934_out0 = v$REGDIN_3350_out0;
assign v$REGDIN_1935_out0 = v$REGDIN_3351_out0;
assign v$MUX5_2882_out0 = v$RET_2207_out0 ? v$REG2_750_out0 : v$MUX4_788_out0;
assign v$MUX5_2883_out0 = v$RET_2208_out0 ? v$REG2_751_out0 : v$MUX4_789_out0;
assign v$NOTUSED_4762_out0 = v$_3346_out1;
assign v$NOTUSED_4763_out0 = v$_3347_out1;
assign v$ControlRequest2_5031_out0 = v$CONTROLREQUEST2_4145_out0;
assign v$_5099_out0 = v$_3126_out1[0:0];
assign v$_5099_out1 = v$_3126_out1[11:11];
assign v$_5100_out0 = v$_3127_out1[0:0];
assign v$_5100_out1 = v$_3127_out1[11:11];
assign v$MUX3_5264_out0 = v$_1569_out0 ? v$MSL_591_out0 : v$IN_2403_out0;
assign v$MUX3_5265_out0 = v$_1570_out0 ? v$MSL_592_out0 : v$IN_2404_out0;
assign v$_1580_out0 = v$ControlRequest2_5031_out0[0:0];
assign v$_1580_out1 = v$ControlRequest2_5031_out0[1:1];
assign v$OUT_1757_out0 = v$MUX1_1435_out0;
assign v$OUT_1758_out0 = v$MUX1_1436_out0;
assign v$_3464_out0 = v$ControlRequest1_214_out0[0:0];
assign v$_3464_out1 = v$ControlRequest1_214_out0[1:1];
assign v$MUX2_3809_out0 = v$_1569_out1 ? v$MUX4_276_out0 : v$MUX3_5264_out0;
assign v$MUX2_3810_out0 = v$_1570_out1 ? v$MUX4_277_out0 : v$MUX3_5265_out0;
assign v$_4723_out0 = v$_5099_out1[0:0];
assign v$_4723_out1 = v$_5099_out1[10:10];
assign v$_4724_out0 = v$_5100_out1[0:0];
assign v$_4724_out1 = v$_5100_out1[10:10];
assign v$RAMADDRMUX_5262_out0 = v$RAMADDRMUX_1479_out0;
assign v$RAMADDRMUX_5263_out0 = v$RAMADDRMUX_1480_out0;
assign v$RAMADDRMUX_613_out0 = v$RAMADDRMUX_5262_out0;
assign v$RAMADDRMUX_614_out0 = v$RAMADDRMUX_5263_out0;
assign v$PRIORITY1_2673_out0 = v$_3464_out1;
assign v$IN_3131_out0 = v$OUT_1757_out0;
assign v$IN_3132_out0 = v$OUT_1758_out0;
assign v$CONTROLREQ1_3719_out0 = v$_3464_out0;
assign v$MUX1_3902_out0 = v$EQ1_1314_out0 ? v$MUX2_3809_out0 : v$IN_2403_out0;
assign v$MUX1_3903_out0 = v$EQ1_1315_out0 ? v$MUX2_3810_out0 : v$IN_2404_out0;
assign v$PRIORITY2_4698_out0 = v$_1580_out1;
assign v$_5048_out0 = v$_4723_out1[0:0];
assign v$_5048_out1 = v$_4723_out1[9:9];
assign v$_5049_out0 = v$_4724_out1[0:0];
assign v$_5049_out1 = v$_4724_out1[9:9];
assign v$CONTROLREQ2_5432_out0 = v$_1580_out0;
assign v$G2_518_out0 = ((v$CONTROLREQ2_5432_out0 && !v$CONTROLREQ1_3719_out0) || (!v$CONTROLREQ2_5432_out0) && v$CONTROLREQ1_3719_out0);
assign v$G1_1258_out0 = v$CONTROLREQ2_5432_out0 && v$CONTROLREQ1_3719_out0;
assign v$_2378_out0 = v$_5048_out1[0:0];
assign v$_2378_out1 = v$_5048_out1[8:8];
assign v$_2379_out0 = v$_5049_out1[0:0];
assign v$_2379_out1 = v$_5049_out1[8:8];
assign v$OUT_3063_out0 = v$MUX1_3902_out0;
assign v$OUT_3064_out0 = v$MUX1_3903_out0;
assign v$RAMADDRMUX_3785_out0 = v$RAMADDRMUX_613_out0;
assign v$RAMADDRMUX_3786_out0 = v$RAMADDRMUX_614_out0;
assign v$IN_4526_out0 = v$IN_3131_out0;
assign v$IN_4527_out0 = v$IN_3132_out0;
assign v$G3_4849_out0 = !((v$PRIORITY1_2673_out0 && !v$PRIORITY2_4698_out0) || (!v$PRIORITY1_2673_out0) && v$PRIORITY2_4698_out0);
assign v$_1080_out0 = v$IN_4526_out0[13:0];
assign v$_1080_out1 = v$IN_4526_out0[15:2];
assign v$_1081_out0 = v$IN_4527_out0[13:0];
assign v$_1081_out1 = v$IN_4527_out0[15:2];
assign v$G4_2999_out0 = v$G3_4849_out0 && v$G1_1258_out0;
assign v$MUX2_3778_out0 = v$G3_4849_out0 ? v$PRIORITYSAME_5355_out0 : v$PRIORITY2_4698_out0;
assign v$MUX1_3966_out0 = v$FETCH_3722_out0 ? v$PC1_987_out0 : v$RAMADDRMUX_3785_out0;
assign v$MUX1_3967_out0 = v$FETCH_3723_out0 ? v$PC1_988_out0 : v$RAMADDRMUX_3786_out0;
assign v$_4250_out0 = v$_2378_out1[0:0];
assign v$_4250_out1 = v$_2378_out1[7:7];
assign v$_4251_out0 = v$_2379_out1[0:0];
assign v$_4251_out1 = v$_2379_out1[7:7];
assign v$_4408_out0 = v$IN_4526_out0[1:0];
assign v$_4408_out1 = v$IN_4526_out0[15:14];
assign v$_4409_out0 = v$IN_4527_out0[1:0];
assign v$_4409_out1 = v$IN_4527_out0[15:14];
assign v$_281_out0 = { v$_4408_out1,v$ZERO_3309_out0 };
assign v$_282_out0 = { v$_4409_out1,v$ZERO_3310_out0 };
assign v$_515_out0 = { v$_4408_out1,v$_4408_out0 };
assign v$_516_out0 = { v$_4409_out1,v$_4409_out0 };
assign v$_1551_out0 = { v$ZERO_3309_out0,v$_1080_out0 };
assign v$_1552_out0 = { v$ZERO_3310_out0,v$_1081_out0 };
assign v$MUX3_2226_out0 = v$G2_518_out0 ? v$CONTROLREQ2_5432_out0 : v$MUX2_3778_out0;
assign v$_2717_out0 = v$_4250_out1[0:0];
assign v$_2717_out1 = v$_4250_out1[6:6];
assign v$_2718_out0 = v$_4251_out1[0:0];
assign v$_2718_out1 = v$_4251_out1[6:6];
assign v$_4457_out0 = v$_1080_out1[0:0];
assign v$_4457_out1 = v$_1080_out1[1:1];
assign v$_4458_out0 = v$_1081_out1[0:0];
assign v$_4458_out1 = v$_1081_out1[1:1];
assign v$PROGRAMADDRESS_4514_out0 = v$MUX1_3966_out0;
assign v$PROGRAMADDRESS_4515_out0 = v$MUX1_3967_out0;
assign v$ROR_1018_out0 = v$_515_out0;
assign v$ROR_1019_out0 = v$_516_out0;
assign v$DM2_1095_out0 = v$MUX3_2226_out0 ? 1'h0 : v$C5_4291_out0;
assign v$DM2_1095_out1 = v$MUX3_2226_out0 ? v$C5_4291_out0 : 1'h0;
assign v$DATAADDRESS_2471_out0 = v$PROGRAMADDRESS_4515_out0;
assign v$DATAADDRESS_2472_out0 = v$PROGRAMADDRESS_4514_out0;
assign v$_2509_out0 = { v$_4457_out1,v$_4457_out1 };
assign v$_2510_out0 = { v$_4458_out1,v$_4458_out1 };
assign v$LSR_3076_out0 = v$_281_out0;
assign v$LSR_3077_out0 = v$_282_out0;
assign v$NA_4715_out0 = v$_4457_out0;
assign v$NA_4716_out0 = v$_4458_out0;
assign v$_5027_out0 = v$_2717_out1[0:0];
assign v$_5027_out1 = v$_2717_out1[5:5];
assign v$_5028_out0 = v$_2718_out1[0:0];
assign v$_5028_out1 = v$_2718_out1[5:5];
assign v$LSL_5349_out0 = v$_1551_out0;
assign v$LSL_5350_out0 = v$_1552_out0;
assign v$_1297_out0 = v$_5027_out1[0:0];
assign v$_1297_out1 = v$_5027_out1[4:4];
assign v$_1298_out0 = v$_5028_out1[0:0];
assign v$_1298_out1 = v$_5028_out1[4:4];
assign v$G7_2850_out0 = v$DM2_1095_out1 && v$CONTROLREQ2_5432_out0;
assign v$_3415_out0 = { v$_4408_out1,v$_2509_out0 };
assign v$_3416_out0 = { v$_4409_out1,v$_2510_out0 };
assign v$G6_4830_out0 = v$CONTROLREQ1_3719_out0 && v$DM2_1095_out0;
assign v$MUX3_4904_out0 = v$_523_out1 ? v$ROR_1018_out0 : v$LSR_3076_out0;
assign v$MUX3_4905_out0 = v$_524_out1 ? v$ROR_1019_out0 : v$LSR_3077_out0;
assign v$_5115_out0 = { v$WRITEDATA_1247_out0,v$DATAADDRESS_2471_out0 };
assign v$_5116_out0 = { v$WRITEDATA_1248_out0,v$DATAADDRESS_2472_out0 };
assign v$CONTROLGRANT1_1722_out0 = v$G6_4830_out0;
assign v$_2654_out0 = { v$_5115_out0,v$WREQUEST_508_out0 };
assign v$_2655_out0 = { v$_5116_out0,v$WREQUEST_509_out0 };
assign v$ASR_2947_out0 = v$_3415_out0;
assign v$ASR_2948_out0 = v$_3416_out0;
assign v$_4804_out0 = v$_1297_out1[0:0];
assign v$_4804_out1 = v$_1297_out1[3:3];
assign v$_4805_out0 = v$_1298_out1[0:0];
assign v$_4805_out1 = v$_1298_out1[3:3];
assign v$CONTROLGRANT2_4822_out0 = v$G7_2850_out0;
assign v$WENDATA_162_out0 = v$_2654_out0;
assign v$WENDATA_163_out0 = v$_2655_out0;
assign v$_223_out0 = v$_4804_out1[0:0];
assign v$_223_out1 = v$_4804_out1[2:2];
assign v$_224_out0 = v$_4805_out1[0:0];
assign v$_224_out1 = v$_4805_out1[2:2];
assign v$CONTROLGRANT2_406_out0 = v$CONTROLGRANT2_4822_out0;
assign v$CONTROLGRANT1_1378_out0 = v$CONTROLGRANT1_1722_out0;
assign v$MUX2_2255_out0 = v$_523_out1 ? v$ASR_2947_out0 : v$LSL_5349_out0;
assign v$MUX2_2256_out0 = v$_524_out1 ? v$ASR_2948_out0 : v$LSL_5350_out0;
assign v$WENDATA1_1446_out0 = v$WENDATA_163_out0;
assign v$_1512_out0 = v$_223_out1[0:0];
assign v$_1512_out1 = v$_223_out1[1:1];
assign v$_1513_out0 = v$_224_out1[0:0];
assign v$_1513_out1 = v$_224_out1[1:1];
assign v$CONTROLGRANT_1832_out0 = v$CONTROLGRANT2_406_out0;
assign v$CONTROLGRANT_1833_out0 = v$CONTROLGRANT1_1378_out0;
assign v$MUX4_1893_out0 = v$_523_out0 ? v$MUX3_4904_out0 : v$MUX2_2255_out0;
assign v$MUX4_1894_out0 = v$_524_out0 ? v$MUX3_4905_out0 : v$MUX2_2256_out0;
assign v$WENDATA2_2308_out0 = v$WENDATA_162_out0;
assign v$WEN$DATA2_3530_out0 = v$WENDATA2_2308_out0;
assign v$WEN$DATA1_3913_out0 = v$WENDATA1_1446_out0;
assign v$DM1_4074_out0 = v$RREQUEST_3720_out0 ? 1'h0 : v$CONTROLGRANT_1832_out0;
assign v$DM1_4074_out1 = v$RREQUEST_3720_out0 ? v$CONTROLGRANT_1832_out0 : 1'h0;
assign v$DM1_4075_out0 = v$RREQUEST_3721_out0 ? 1'h0 : v$CONTROLGRANT_1833_out0;
assign v$DM1_4075_out1 = v$RREQUEST_3721_out0 ? v$CONTROLGRANT_1833_out0 : 1'h0;
assign v$MUX1_4868_out0 = v$EN_1424_out0 ? v$MUX4_1893_out0 : v$IN_4526_out0;
assign v$MUX1_4869_out0 = v$EN_1425_out0 ? v$MUX4_1894_out0 : v$IN_4527_out0;
assign v$WRITECOMPLETE_203_out0 = v$DM1_4074_out0;
assign v$WRITECOMPLETE_204_out0 = v$DM1_4075_out0;
assign v$OUT_1077_out0 = v$MUX1_4868_out0;
assign v$OUT_1078_out0 = v$MUX1_4869_out0;
assign v$CONTROLPROTOCAL2_1243_out0 = v$WEN$DATA2_3530_out0;
assign v$READVALID_2915_out0 = v$DM1_4074_out1;
assign v$READVALID_2916_out0 = v$DM1_4075_out1;
assign v$CONTROLPROTOCAL1_4086_out0 = v$WEN$DATA1_3913_out0;
assign v$READVALID_178_out0 = v$READVALID_2916_out0;
assign v$READVALID_179_out0 = v$READVALID_2915_out0;
assign v$WRITECOMPLETE_487_out0 = v$WRITECOMPLETE_204_out0;
assign v$WRITECOMPLETE_488_out0 = v$WRITECOMPLETE_203_out0;
assign v$MUX1_2742_out0 = v$MUX3_2226_out0 ? v$CONTROLPROTOCAL2_1243_out0 : v$CONTROLPROTOCAL1_4086_out0;
assign v$IN_4914_out0 = v$OUT_1077_out0;
assign v$IN_4915_out0 = v$OUT_1078_out0;
assign v$IN_353_out0 = v$IN_4914_out0;
assign v$IN_354_out0 = v$IN_4915_out0;
assign v$_3365_out0 = v$MUX1_2742_out0[27:0];
assign v$_3365_out1 = v$MUX1_2742_out0[28:1];
assign v$G11_4253_out0 = ((v$READVALID_178_out0 && !v$READREQ_2930_out0) || (!v$READVALID_178_out0) && v$READREQ_2930_out0);
assign v$G11_4254_out0 = ((v$READVALID_179_out0 && !v$READREQ_2931_out0) || (!v$READVALID_179_out0) && v$READREQ_2931_out0);
assign v$G12_5211_out0 = ((v$WRITEREQ_2132_out0 && !v$WRITECOMPLETE_487_out0) || (!v$WRITEREQ_2132_out0) && v$WRITECOMPLETE_487_out0);
assign v$G12_5212_out0 = ((v$WRITEREQ_2133_out0 && !v$WRITECOMPLETE_488_out0) || (!v$WRITEREQ_2133_out0) && v$WRITECOMPLETE_488_out0);
assign v$G13_326_out0 = v$G11_4253_out0 || v$G12_5211_out0;
assign v$G13_327_out0 = v$G11_4254_out0 || v$G12_5212_out0;
assign v$_1236_out0 = v$_3365_out0[15:0];
assign v$_1236_out1 = v$_3365_out0[27:12];
assign v$_2787_out0 = v$IN_353_out0[3:0];
assign v$_2787_out1 = v$IN_353_out0[15:12];
assign v$_2788_out0 = v$IN_354_out0[3:0];
assign v$_2788_out1 = v$IN_354_out0[15:12];
assign v$WRITEENABLE_3250_out0 = v$_3365_out1;
assign v$_3422_out0 = v$IN_353_out0[11:0];
assign v$_3422_out1 = v$IN_353_out0[15:4];
assign v$_3423_out0 = v$IN_354_out0[11:0];
assign v$_3423_out1 = v$IN_354_out0[15:4];
assign v$_636_out0 = { v$ZERO_3207_out0,v$_3422_out0 };
assign v$_637_out0 = { v$ZERO_3208_out0,v$_3423_out0 };
assign v$WRITEENABLE_790_out0 = v$WRITEENABLE_3250_out0;
assign v$WRITEDATA_813_out0 = v$_1236_out0;
assign v$ADDRESS_1313_out0 = v$_1236_out1;
assign v$_4151_out0 = { v$_2787_out1,v$_2787_out0 };
assign v$_4152_out0 = { v$_2788_out1,v$_2788_out0 };
assign v$_4153_out0 = { v$_2787_out1,v$ZERO_3207_out0 };
assign v$_4154_out0 = { v$_2788_out1,v$ZERO_3208_out0 };
assign v$_5062_out0 = v$_3422_out1[2:0];
assign v$_5062_out1 = v$_3422_out1[3:1];
assign v$_5063_out0 = v$_3423_out1[2:0];
assign v$_5063_out1 = v$_3423_out1[3:1];
assign v$STALL_5393_out0 = v$G13_326_out0;
assign v$STALL_5394_out0 = v$G13_327_out0;
assign v$WRITEDATA_1328_out0 = v$WRITEDATA_813_out0;
assign v$DMADDRESS_1885_out0 = v$ADDRESS_1313_out0;
assign v$LSL_2051_out0 = v$_636_out0;
assign v$LSL_2052_out0 = v$_637_out0;
assign v$STALL_2382_out0 = v$STALL_5393_out0;
assign v$STALL_2383_out0 = v$STALL_5394_out0;
assign v$_2476_out0 = { v$_5062_out1,v$_5062_out1 };
assign v$_2477_out0 = { v$_5063_out1,v$_5063_out1 };
assign v$ROR_2513_out0 = v$_4151_out0;
assign v$ROR_2514_out0 = v$_4152_out0;
assign v$LSR_2641_out0 = v$_4153_out0;
assign v$LSR_2642_out0 = v$_4154_out0;
assign v$STALL_2680_out0 = v$STALL_5393_out0;
assign v$STALL_2681_out0 = v$STALL_5394_out0;
assign v$NA_3557_out0 = v$_5062_out0;
assign v$NA_3558_out0 = v$_5063_out0;
assign v$STALL_3987_out0 = v$STALL_5393_out0;
assign v$STALL_3988_out0 = v$STALL_5394_out0;
assign v$STALL_4418_out0 = v$STALL_5393_out0;
assign v$STALL_4419_out0 = v$STALL_5394_out0;
assign v$STALL_4480_out0 = v$STALL_5393_out0;
assign v$STALL_4481_out0 = v$STALL_5394_out0;
assign v$ADDRESS_4_out0 = v$DMADDRESS_1885_out0;
assign v$_1527_out0 = { v$_2476_out0,v$_2476_out0 };
assign v$_1528_out0 = { v$_2477_out0,v$_2477_out0 };
assign v$WDATA_1785_out0 = v$WRITEDATA_1328_out0;
assign v$MUX3_2384_out0 = v$_1244_out1 ? v$ROR_2513_out0 : v$LSR_2641_out0;
assign v$MUX3_2385_out0 = v$_1245_out1 ? v$ROR_2514_out0 : v$LSR_2642_out0;
assign v$STALL2_2936_out0 = v$STALL_2681_out0;
assign v$STALL1_3563_out0 = v$STALL_2680_out0;
assign v$G9_4580_out0 = ! v$STALL_4418_out0;
assign v$G9_4581_out0 = ! v$STALL_4419_out0;
assign v$STALL_4645_out0 = v$STALL_4480_out0;
assign v$STALL_4646_out0 = v$STALL_4481_out0;
assign v$STALL_5064_out0 = v$STALL_3987_out0;
assign v$STALL_5065_out0 = v$STALL_3988_out0;
assign v$_956_out0 = { v$_2787_out1,v$_1527_out0 };
assign v$_957_out0 = { v$_2788_out1,v$_1528_out0 };
assign v$MUX5_2340_out0 = v$STALL_5064_out0 ? v$G1_909_out0 : v$C1_4332_out0;
assign v$MUX5_2341_out0 = v$STALL_5065_out0 ? v$G1_910_out0 : v$C1_4333_out0;
assign v$MUX2_2396_out0 = v$STALL_5064_out0 ? v$C1_4332_out0 : v$G1_909_out0;
assign v$MUX2_2397_out0 = v$STALL_5065_out0 ? v$C1_4333_out0 : v$G1_910_out0;
assign v$MUX7_2479_out0 = v$STALL_5064_out0 ? v$_1749_out0 : v$C1_4332_out0;
assign v$MUX7_2480_out0 = v$STALL_5065_out0 ? v$_1750_out0 : v$C1_4333_out0;
assign v$MUX8_2951_out0 = v$STALL_5064_out0 ? v$C1_4332_out0 : v$G1_909_out0;
assign v$MUX8_2952_out0 = v$STALL_5065_out0 ? v$C1_4333_out0 : v$G1_910_out0;
assign v$G10_3240_out0 = v$EXEC2_3776_out0 && v$G9_4580_out0;
assign v$G10_3241_out0 = v$EXEC2_3777_out0 && v$G9_4581_out0;
assign v$WDATA_4407_out0 = v$WDATA_1785_out0;
assign v$ADDRESS_4829_out0 = v$ADDRESS_4_out0;
assign v$ASR_232_out0 = v$_956_out0;
assign v$ASR_233_out0 = v$_957_out0;
assign v$ADDRESS_2096_out0 = v$ADDRESS_4829_out0;
assign v$MUX6_2954_out0 = v$_4077_out0 ? v$MUX5_2340_out0 : v$MUX8_2951_out0;
assign v$MUX6_2955_out0 = v$_4078_out0 ? v$MUX5_2341_out0 : v$MUX8_2952_out0;
assign v$MUX3_3424_out0 = v$_4077_out0 ? v$MUX2_2396_out0 : v$MUX7_2479_out0;
assign v$MUX3_3425_out0 = v$_4078_out0 ? v$MUX2_2397_out0 : v$MUX7_2480_out0;
assign v$EQ3_415_out0 = v$ADDRESS_2096_out0 == 12'h902;
assign v$EQ5_694_out0 = v$ADDRESS_2096_out0 == 12'h904;
assign v$EQ4_3762_out0 = v$ADDRESS_2096_out0 == 12'h903;
assign v$_4258_out0 = { v$MUX6_2954_out0,v$MUX3_3424_out0 };
assign v$_4259_out0 = { v$MUX6_2955_out0,v$MUX3_3425_out0 };
assign v$MUX2_4708_out0 = v$_1244_out1 ? v$ASR_232_out0 : v$LSL_2051_out0;
assign v$MUX2_4709_out0 = v$_1245_out1 ? v$ASR_233_out0 : v$LSL_2052_out0;
assign v$EQ1_4874_out0 = v$ADDRESS_2096_out0 == 12'h900;
assign v$EQ2_5208_out0 = v$ADDRESS_2096_out0 == 12'h901;
assign v$MUX4_1067_out0 = v$_1244_out0 ? v$MUX3_2384_out0 : v$MUX2_4708_out0;
assign v$MUX4_1068_out0 = v$_1245_out0 ? v$MUX3_2385_out0 : v$MUX2_4709_out0;
assign v$LOAD_2672_out0 = v$EQ5_694_out0;
assign v$ADDB_3280_out0 = v$EQ2_5208_out0;
assign v$MULTB_3304_out0 = v$EQ4_3762_out0;
assign v$A_3523_out0 = v$EQ1_4874_out0;
assign v$Q1_4523_out0 = v$_4258_out0;
assign v$Q1_4524_out0 = v$_4259_out0;
assign v$SUBB_4737_out0 = v$EQ3_415_out0;
assign v$G13_254_out0 = v$FF1_5073_out0 || v$SUBB_4737_out0;
assign v$G15_1113_out0 = v$A_3523_out0 && v$CYC1_3443_out0;
assign v$G3_1413_out0 = v$ADDB_3280_out0 || v$SUBB_4737_out0;
assign v$LOAD_1490_out0 = v$LOAD_2672_out0;
assign v$A_2566_out0 = v$A_3523_out0;
assign v$G14_2733_out0 = v$FF2_3403_out0 || v$MULTB_3304_out0;
assign v$D_5138_out0 = v$Q1_4523_out0;
assign v$D_5139_out0 = v$Q1_4524_out0;
assign v$MUX1_5298_out0 = v$EN_4955_out0 ? v$MUX4_1067_out0 : v$IN_353_out0;
assign v$MUX1_5299_out0 = v$EN_4956_out0 ? v$MUX4_1068_out0 : v$IN_354_out0;
assign v$SUB_510_out0 = v$G13_254_out0;
assign v$MULT_991_out0 = v$G14_2733_out0;
assign v$G8_1311_out0 = v$CYC2_1461_out0 || v$G15_1113_out0;
assign v$A_2182_out0 = v$A_2566_out0;
assign v$_4344_out0 = v$D_5138_out0[0:0];
assign v$_4344_out1 = v$D_5138_out0[1:1];
assign v$_4345_out0 = v$D_5139_out0[0:0];
assign v$_4345_out1 = v$D_5139_out0[1:1];
assign v$G4_5249_out0 = ! v$A_2566_out0;
assign v$OUT_5294_out0 = v$MUX1_5298_out0;
assign v$OUT_5295_out0 = v$MUX1_5299_out0;
assign v$G4_5336_out0 = v$G3_1413_out0 || v$MULTB_3304_out0;
assign v$DM1_492_out0 = v$MULT_991_out0 ? 16'h0 : v$REG1_1106_out0;
assign v$DM1_492_out1 = v$MULT_991_out0 ? v$REG1_1106_out0 : 16'h0;
assign v$NA_1199_out0 = v$G4_5249_out0;
assign v$MULT_1828_out0 = v$MULT_991_out0;
assign v$SUBTRACTOR_3177_out0 = v$SUB_510_out0;
assign v$DM2_3561_out0 = v$MULT_991_out0 ? 16'h0 : v$REG2_5309_out0;
assign v$DM2_3561_out1 = v$MULT_991_out0 ? v$REG2_5309_out0 : 16'h0;
assign v$IN_4576_out0 = v$OUT_5294_out0;
assign v$IN_4577_out0 = v$OUT_5295_out0;
assign v$B_4780_out0 = v$G4_5336_out0;
assign v$SUB_5242_out0 = v$SUB_510_out0;
assign v$MULT_49_out0 = v$MULT_1828_out0;
assign v$B_147_out0 = v$B_4780_out0;
assign v$A_602_out0 = v$DM1_492_out1;
assign v$A_749_out0 = v$DM1_492_out0;
assign v$G16_971_out0 = v$B_4780_out0 && v$CYC1_3443_out0;
assign v$IN_1026_out0 = v$IN_4576_out0;
assign v$IN_1027_out0 = v$IN_4577_out0;
assign v$SUBTRACTOR_1459_out0 = v$SUBTRACTOR_3177_out0;
assign v$B_2005_out0 = v$DM2_3561_out1;
assign v$SUB_3499_out0 = v$SUB_5242_out0;
assign v$G15_4791_out0 = v$NQ0_5_out0 && v$NA_1199_out0;
assign v$B_5337_out0 = v$DM2_3561_out0;
assign v$G5_1623_out0 = ! v$B_147_out0;
assign v$A_2331_out0 = v$A_749_out0;
assign v$_3006_out0 = v$IN_1026_out0[7:0];
assign v$_3006_out1 = v$IN_1026_out0[15:8];
assign v$_3007_out0 = v$IN_1027_out0[7:0];
assign v$_3007_out1 = v$IN_1027_out0[15:8];
assign v$B_3539_out0 = v$B_5337_out0;
assign v$B_3975_out0 = v$B_147_out0;
assign v$B_5057_out0 = v$B_2005_out0;
assign v$A_5334_out0 = v$A_602_out0;
assign v$NB_547_out0 = v$G5_1623_out0;
assign v$SEL2_814_out0 = v$B_3539_out0[14:10];
assign v$SEL2_970_out0 = v$B_3539_out0[9:0];
assign v$SEL1_1118_out0 = v$B_5057_out0[14:10];
assign v$SEL4_1457_out0 = v$A_5334_out0[14:10];
assign v$G16_2159_out0 = v$G15_4791_out0 && v$B_3975_out0;
assign v$SEL1_2457_out0 = v$A_2331_out0[9:0];
assign v$SEL2_2921_out0 = v$B_5057_out0[9:0];
assign v$SEL3_3116_out0 = v$A_5334_out0[9:0];
assign v$7TO0_3572_out0 = v$_3006_out0;
assign v$7TO0_3573_out0 = v$_3007_out0;
assign v$SEL1_3647_out0 = v$A_2331_out0[14:10];
assign v$SEL6_3676_out0 = v$B_5057_out0[15:15];
assign v$SEL5_3993_out0 = v$A_5334_out0[15:15];
assign v$SEL1_4138_out0 = v$A_2331_out0[15:15];
assign v$15TO8_5054_out0 = v$_3006_out1;
assign v$15TO8_5055_out0 = v$_3007_out1;
assign v$SEL2_5321_out0 = v$B_3539_out0[15:15];
assign v$_377_out0 = { v$ZERO_295_out0,v$7TO0_3572_out0 };
assign v$_378_out0 = { v$ZERO_296_out0,v$7TO0_3573_out0 };
assign v$EXPA_1502_out0 = v$SEL4_1457_out0;
assign v$FRACA_1548_out0 = v$SEL1_2457_out0;
assign v$FRACA_1732_out0 = v$SEL3_3116_out0;
assign v$SGNB_1810_out0 = v$SEL2_5321_out0;
assign v$Q$_2632_out0 = v$G16_2159_out0;
assign v$EXPB_3248_out0 = v$SEL2_814_out0;
assign v$_3447_out0 = { v$15TO8_5054_out0,v$ZERO_295_out0 };
assign v$_3448_out0 = { v$15TO8_5055_out0,v$ZERO_296_out0 };
assign v$FRACB_3484_out0 = v$SEL2_2921_out0;
assign v$SGNB_3492_out0 = v$SEL6_3676_out0;
assign v$_3641_out0 = { v$15TO8_5054_out0,v$7TO0_3572_out0 };
assign v$_3642_out0 = { v$15TO8_5055_out0,v$7TO0_3573_out0 };
assign v$FRACB_3827_out0 = v$SEL2_970_out0;
assign v$_3832_out0 = v$15TO8_5054_out0[6:0];
assign v$_3832_out1 = v$15TO8_5054_out0[7:1];
assign v$_3833_out0 = v$15TO8_5055_out0[6:0];
assign v$_3833_out1 = v$15TO8_5055_out0[7:1];
assign v$EXPB_3876_out0 = v$SEL1_1118_out0;
assign v$SGNA_3917_out0 = v$SEL5_3993_out0;
assign v$SGNA_4123_out0 = v$SEL1_4138_out0;
assign v$EXPA_4353_out0 = v$SEL1_3647_out0;
assign v$XOR1_679_out0 = v$SGNA_4123_out0 ^ v$SGNB_1810_out0;
assign v$_1050_out0 = { v$_3832_out1,v$_3832_out1 };
assign v$_1051_out0 = { v$_3833_out1,v$_3833_out1 };
assign v$EXPOA_1226_out0 = v$EXPA_1502_out0;
assign v$G2_1242_out0 = ((v$SGNA_3917_out0 && !v$SGNB_3492_out0) || (!v$SGNA_3917_out0) && v$SGNB_3492_out0);
assign v$LSL_1395_out0 = v$_377_out0;
assign v$LSL_1396_out0 = v$_378_out0;
assign v$EXPOB_1579_out0 = v$EXPB_3876_out0;
assign v$NA_1621_out0 = v$_3832_out0;
assign v$NA_1622_out0 = v$_3833_out0;
assign v$EXPOA_2078_out0 = v$EXPA_4353_out0;
assign v$LSR_2177_out0 = v$_3447_out0;
assign v$LSR_2178_out0 = v$_3448_out0;
assign v$ROR_2757_out0 = v$_3641_out0;
assign v$ROR_2758_out0 = v$_3642_out0;
assign v$EXPOB_5159_out0 = v$EXPB_3248_out0;
assign v$EQ6_612_out0 = v$EXPOB_1579_out0 == 5'h0;
assign v$G1_795_out0 = ! v$XOR1_679_out0;
assign v$EXPONENTA_1574_out0 = v$EXPOA_2078_out0;
assign v$EQ7_1762_out0 = v$EXPOA_1226_out0 == 5'h0;
assign v$EXPOA_1813_out0 = v$EXPOA_1226_out0;
assign v$EXPONENTB_2080_out0 = v$EXPOB_5159_out0;
assign v$_2328_out0 = { v$_1050_out0,v$_1050_out0 };
assign v$_2329_out0 = { v$_1051_out0,v$_1051_out0 };
assign v$SGNOUT_2961_out0 = v$XOR1_679_out0;
assign v$EQ2_3018_out0 = v$EXPOB_1579_out0 == 5'h1f;
assign v$MUX3_3205_out0 = v$_2186_out1 ? v$ROR_2757_out0 : v$LSR_2177_out0;
assign v$MUX3_3206_out0 = v$_2187_out1 ? v$ROR_2758_out0 : v$LSR_2178_out0;
assign v$SUB_3371_out0 = v$XOR1_679_out0;
assign v$EXPOB_3402_out0 = v$EXPOB_1579_out0;
assign v$SGN_3620_out0 = v$G2_1242_out0;
assign v$EQ1_5213_out0 = v$EXPOA_1226_out0 == 5'h1f;
assign v$_14_out0 = { v$_2328_out0,v$_2328_out0 };
assign v$_15_out0 = { v$_2329_out0,v$_2329_out0 };
assign v$ADD_497_out0 = v$G1_795_out0;
assign v$INFINITYB_1517_out0 = v$EQ2_3018_out0;
assign v$EQ9_2267_out0 = v$EXPONENTB_2080_out0 == 5'h0;
assign v$MUX3_2558_out0 = v$EQ6_612_out0 ? v$C9_1415_out0 : v$EXPOB_1579_out0;
assign v$INFINITYA_2940_out0 = v$EQ1_5213_out0;
assign v$EQ3_3053_out0 = v$EXPONENTA_1574_out0 == 5'h0;
assign v$EQ8_3303_out0 = v$EXPONENTA_1574_out0 == 5'h0;
assign v$SIGNOPERATION_3729_out0 = v$SGNOUT_2961_out0;
assign v$EQ4_3781_out0 = v$EXPONENTA_1574_out0 == 5'h1f;
assign v$EQ5_3879_out0 = v$EXPOB_3402_out0 == 5'h0;
assign v$EQ3_4431_out0 = v$EXPOA_1813_out0 == 5'h0;
assign v$EQ6_4710_out0 = v$EXPONENTB_2080_out0 == 5'h0;
assign v$EQ5_4729_out0 = v$EXPONENTB_2080_out0 == 5'h1f;
assign v$MUX4_4779_out0 = v$EQ7_1762_out0 ? v$C10_2986_out0 : v$EXPOA_1226_out0;
assign v$ZERO_778_out0 = v$EQ3_3053_out0;
assign v$G4_1418_out0 = ((v$SUBTRACTOR_1459_out0 && !v$SIGNOPERATION_3729_out0) || (!v$SUBTRACTOR_1459_out0) && v$SIGNOPERATION_3729_out0);
assign v$ADDONEA_1550_out0 = v$EQ8_3303_out0;
assign v$INFINITY16_2098_out0 = v$EQ5_4729_out0;
assign v$ZERO_2473_out0 = v$EQ3_4431_out0;
assign v$ADDONEB_2625_out0 = v$EQ9_2267_out0;
assign v$_3061_out0 = { v$15TO8_5054_out0,v$_14_out0 };
assign v$_3062_out0 = { v$15TO8_5055_out0,v$_15_out0 };
assign v$ZERO14_3688_out0 = v$EQ5_3879_out0;
assign v$INFINITY_4150_out0 = v$EQ4_3781_out0;
assign v$ZERO14_4652_out0 = v$EQ6_4710_out0;
assign v$G1_5051_out0 = v$INFINITYA_2940_out0 || v$INFINITYB_1517_out0;
assign {v$A1_5395_out1,v$A1_5395_out0 } = v$MUX4_4779_out0 + v$MUX3_2558_out0 + v$C1_1360_out0;
assign v$_482_out0 = { v$A1_5395_out0,v$A1_5395_out1 };
assign v$G1_695_out0 = ! v$ZERO_778_out0;
assign v$G2_763_out0 = ! v$ZERO14_3688_out0;
assign v$ASR_834_out0 = v$_3061_out0;
assign v$ASR_835_out0 = v$_3062_out0;
assign v$INFINITY_1025_out0 = v$G1_5051_out0;
assign v$MUX5_1030_out0 = v$ADDONEB_2625_out0 ? v$C9_3886_out0 : v$EXPONENTB_2080_out0;
assign v$MUX4_1182_out0 = v$ADDONEA_1550_out0 ? v$C9_3886_out0 : v$EXPONENTA_1574_out0;
assign v$INFINITY_2028_out0 = v$INFINITY_4150_out0;
assign v$G1_3986_out0 = ! v$ZERO_2473_out0;
assign v$INFINITY2_4485_out0 = v$INFINITY16_2098_out0;
assign v$SUB_4899_out0 = v$G4_1418_out0;
assign v$G2_5400_out0 = ! v$ZERO14_4652_out0;
assign v$XOR1_16_out0 = v$C1_2374_out0 ^ v$MUX5_1030_out0;
assign v$MUX2_155_out0 = v$G2_5400_out0 ? v$C4_1000_out0 : v$C5_4435_out0;
assign v$INFINITY_231_out0 = v$INFINITY_2028_out0;
assign v$MUX2_792_out0 = v$_2186_out1 ? v$ASR_834_out0 : v$LSL_1395_out0;
assign v$MUX2_793_out0 = v$_2187_out1 ? v$ASR_835_out0 : v$LSL_1396_out0;
assign v$MUX2_843_out0 = v$G1_3986_out0 ? v$C7_4222_out0 : v$C6_297_out0;
assign v$INFINITYB_1096_out0 = v$INFINITY2_4485_out0;
assign v$_1127_out0 = { v$_482_out0,v$C4_2185_out0 };
assign v$MUX1_3538_out0 = v$G2_763_out0 ? v$C5_4513_out0 : v$C8_1437_out0;
assign v$MUX1_3730_out0 = v$G1_695_out0 ? v$C3_3579_out0 : v$C2_1970_out0;
assign v$MUX1_4000_out0 = v$SUB_4899_out0 ? v$C1_4937_out0 : v$C2_743_out0;
assign v$G2_4803_out0 = ! v$SUB_4899_out0;
assign v$FRACTIONINTA_348_out0 = v$MUX2_843_out0;
assign v$FRACTIONINTA_631_out0 = v$MUX1_3730_out0;
assign v$G1_706_out0 = v$INFINITY_231_out0 || v$INFINITYB_1096_out0;
assign v$MUX4_1306_out0 = v$_2186_out0 ? v$MUX3_3205_out0 : v$MUX2_792_out0;
assign v$MUX4_1307_out0 = v$_2187_out0 ? v$MUX3_3206_out0 : v$MUX2_793_out0;
assign v$FRACTIONINTB_1578_out0 = v$MUX1_3538_out0;
assign v$FRACTIONINTB_3004_out0 = v$MUX2_155_out0;
assign {v$comparator_4432_out1,v$comparator_4432_out0 } = v$MUX4_1182_out0 + v$XOR1_16_out0 + v$C0_2686_out0;
assign {v$A2_4445_out1,v$A2_4445_out0 } = v$_1127_out0 + v$C2_4547_out0 + v$C3_3433_out0;
assign v$X1_165_out0 = v$A2_4445_out1;
assign v$_811_out0 = { v$FRACB_3827_out0,v$FRACTIONINTB_3004_out0 };
assign v$EQ7_1017_out0 = v$comparator_4432_out0 == 5'h0;
assign v$G5_2063_out0 = v$FRACTIONINTA_348_out0 && v$FRACTIONINTB_1578_out0;
assign v$_2070_out0 = { v$FRACB_3484_out0,v$FRACTIONINTB_1578_out0 };
assign v$EXPONENTDIFFERENCE13_2330_out0 = v$comparator_4432_out0;
assign v$EXPO_2336_out0 = v$A2_4445_out0;
assign v$EQ1_2759_out0 = v$comparator_4432_out1 == 1'h0;
assign v$_3051_out0 = { v$FRACA_1548_out0,v$FRACTIONINTA_631_out0 };
assign v$_3831_out0 = { v$FRACA_1732_out0,v$FRACTIONINTA_348_out0 };
assign v$EQ0_4033_out0 = v$comparator_4432_out1 == 1'h1;
assign v$MUX1_4389_out0 = v$EN_5416_out0 ? v$MUX4_1306_out0 : v$IN_1026_out0;
assign v$MUX1_4390_out0 = v$EN_5417_out0 ? v$MUX4_1307_out0 : v$IN_1027_out0;
assign v$EQ2_5209_out0 = v$comparator_4432_out0 == 5'h0;
assign v$EXPO_44_out0 = v$EXPO_2336_out0;
assign v$FRAC11A_154_out0 = v$_3051_out0;
assign v$MULTIPLIER_1024_out0 = v$_2070_out0;
assign v$G3_1542_out0 = ! v$EQ7_1017_out0;
assign {v$A1_1910_out1,v$A1_1910_out0 } = v$EXPONENTDIFFERENCE13_2330_out0 + v$C7_2066_out0 + v$C8_4120_out0;
assign v$ABEQUAL_2065_out0 = v$EQ2_5209_out0;
assign v$FRAC11B_2912_out0 = v$_811_out0;
assign v$G6_4376_out0 = ! v$G5_2063_out0;
assign v$ASMALLER_4525_out0 = v$EQ1_2759_out0;
assign v$OUT_4569_out0 = v$MUX1_4389_out0;
assign v$OUT_4570_out0 = v$MUX1_4390_out0;
assign v$MULTIPLICAND_5224_out0 = v$_3831_out0;
assign v$$EXPONENT_225_out0 = v$EXPO_44_out0;
assign v$ABEQUAL_341_out0 = v$ABEQUAL_2065_out0;
assign v$G4_615_out0 = v$EQ0_4033_out0 && v$G3_1542_out0;
assign v$X_1667_out0 = v$A1_1910_out1;
assign v$MUX2_2169_out0 = v$EQ1_3645_out0 ? v$OUT_3063_out0 : v$OUT_4569_out0;
assign v$MUX2_2170_out0 = v$EQ1_3646_out0 ? v$OUT_3064_out0 : v$OUT_4570_out0;
assign v$MULTISHIFT_2679_out0 = v$G6_4376_out0;
assign v$_3936_out0 = { v$SGNA_4123_out0,v$FRAC11A_154_out0 };
assign v$FRACB_4130_out0 = v$MULTIPLIER_1024_out0;
assign v$XOR2_4394_out0 = v$C1_1312_out0 ^ v$FRAC11B_2912_out0;
assign v$ASMALLER_4819_out0 = v$ASMALLER_4525_out0;
assign v$FRACA_4929_out0 = v$MULTIPLICAND_5224_out0;
assign v$_4930_out0 = { v$SGNB_1810_out0,v$FRAC11B_2912_out0 };
assign v$XOR2_5112_out0 = v$C6_3481_out0 ^ v$A1_1910_out0;
assign v$EXPONENT_5290_out0 = v$EXPO_44_out0;
assign v$EXPONENT_5297_out0 = v$EXPO_44_out0;
assign v$SEL4_676_out0 = v$EXPONENT_5297_out0[5:0];
assign v$SEL1_744_out0 = v$$EXPONENT_225_out0[6:6];
assign v$B_951_out0 = v$FRACB_4130_out0;
assign v$XOR1_1741_out0 = v$$EXPONENT_225_out0 ^ v$C13_1573_out0;
assign v$SHIFTOUT_1795_out0 = v$MUX2_2169_out0;
assign v$SHIFTOUT_1796_out0 = v$MUX2_2170_out0;
assign v$A_1802_out0 = v$FRACA_4929_out0;
assign v$ASMALLER_2055_out0 = v$ASMALLER_4819_out0;
assign {v$A1_4358_out1,v$A1_4358_out0 } = v$FRAC11A_154_out0 + v$XOR2_4394_out0 + v$C0_4802_out0;
assign v$ABIGGER_4757_out0 = v$G4_615_out0;
assign v$EXPONENT_5089_out0 = v$EXPONENT_5290_out0;
assign v$SEL3_5279_out0 = v$EXPONENT_5297_out0[6:6];
assign v$X_3_out0 = v$A1_4358_out0;
assign v$SEL7_105_out0 = v$B_951_out0[10:10];
assign v$SEL6_227_out0 = v$B_951_out0[5:5];
assign v$A_470_out0 = v$A_1802_out0;
assign v$A_471_out0 = v$A_1802_out0;
assign v$A_472_out0 = v$A_1802_out0;
assign v$A_473_out0 = v$A_1802_out0;
assign v$A_474_out0 = v$A_1802_out0;
assign v$A_475_out0 = v$A_1802_out0;
assign v$A_476_out0 = v$A_1802_out0;
assign v$A_477_out0 = v$A_1802_out0;
assign v$A_478_out0 = v$A_1802_out0;
assign v$A_479_out0 = v$A_1802_out0;
assign v$A_480_out0 = v$A_1802_out0;
assign v$MUX3_527_out0 = v$ASMALLER_2055_out0 ? v$EXPB_3248_out0 : v$EXPA_4353_out0;
assign v$EQ1_1321_out0 = v$A1_4358_out1 == 1'h0;
assign v$SEL11_1602_out0 = v$B_951_out0[7:7];
assign v$_2023_out0 = { v$EXPONENT_5089_out0,v$C19_4917_out0 };
assign {v$A1_2039_out1,v$A1_2039_out0 } = v$XOR1_1741_out0 + v$C15_4273_out0 + v$C14_3974_out0;
assign v$SEL4_2184_out0 = v$B_951_out0[3:3];
assign v$ABIGGER_2412_out0 = v$ABIGGER_4757_out0;
assign v$OP2_2722_out0 = v$SHIFTOUT_1795_out0;
assign v$OP2_2723_out0 = v$SHIFTOUT_1796_out0;
assign v$SEL1_3332_out0 = v$B_951_out0[0:0];
assign v$SEL8_3411_out0 = v$B_951_out0[8:8];
assign v$NONVALID_3848_out0 = v$SEL3_5279_out0;
assign v$SEL9_3961_out0 = v$B_951_out0[6:6];
assign v$SEL2_3962_out0 = v$B_951_out0[1:1];
assign v$MUX3_4060_out0 = v$ABIGGER_4757_out0 ? v$EXPONENTDIFFERENCE13_2330_out0 : v$XOR2_5112_out0;
assign v$SEL5_4204_out0 = v$B_951_out0[4:4];
assign v$SEL3_4260_out0 = v$B_951_out0[2:2];
assign v$SEL10_4314_out0 = v$B_951_out0[9:9];
assign v$NEGATIVEMODE_5050_out0 = v$SEL1_744_out0;
assign v$NEGATIVEMODE_394_out0 = v$NEGATIVEMODE_5050_out0;
assign v$ABSOLUTE_486_out0 = v$A1_2039_out0;
assign v$_1265_out0 = v$A_470_out0[0:0];
assign v$_1265_out1 = v$A_470_out0[10:10];
assign v$_1266_out0 = v$A_471_out0[0:0];
assign v$_1266_out1 = v$A_471_out0[10:10];
assign v$_1267_out0 = v$A_472_out0[0:0];
assign v$_1267_out1 = v$A_472_out0[10:10];
assign v$_1268_out0 = v$A_473_out0[0:0];
assign v$_1268_out1 = v$A_473_out0[10:10];
assign v$_1269_out0 = v$A_474_out0[0:0];
assign v$_1269_out1 = v$A_474_out0[10:10];
assign v$_1270_out0 = v$A_475_out0[0:0];
assign v$_1270_out1 = v$A_475_out0[10:10];
assign v$_1271_out0 = v$A_476_out0[0:0];
assign v$_1271_out1 = v$A_476_out0[10:10];
assign v$_1272_out0 = v$A_477_out0[0:0];
assign v$_1272_out1 = v$A_477_out0[10:10];
assign v$_1273_out0 = v$A_478_out0[0:0];
assign v$_1273_out1 = v$A_478_out0[10:10];
assign v$_1274_out0 = v$A_479_out0[0:0];
assign v$_1274_out1 = v$A_479_out0[10:10];
assign v$_1275_out0 = v$A_480_out0[0:0];
assign v$_1275_out1 = v$A_480_out0[10:10];
assign v$NONVALID_1544_out0 = v$NONVALID_3848_out0;
assign v$BIGGEREXPO_1814_out0 = v$MUX3_527_out0;
assign v$NOTUSE_2079_out0 = v$A1_2039_out1;
assign v$Asmaller_2247_out0 = v$EQ1_1321_out0;
assign v$OP2_2995_out0 = v$OP2_2722_out0;
assign v$OP2_2996_out0 = v$OP2_2723_out0;
assign v$B_3507_out0 = v$SEL11_1602_out0;
assign v$B_3508_out0 = v$SEL1_3332_out0;
assign v$B_3509_out0 = v$SEL2_3962_out0;
assign v$B_3510_out0 = v$SEL3_4260_out0;
assign v$B_3511_out0 = v$SEL9_3961_out0;
assign v$B_3512_out0 = v$SEL10_4314_out0;
assign v$B_3513_out0 = v$SEL4_2184_out0;
assign v$B_3514_out0 = v$SEL7_105_out0;
assign v$B_3515_out0 = v$SEL5_4204_out0;
assign v$B_3516_out0 = v$SEL8_3411_out0;
assign v$B_3517_out0 = v$SEL6_227_out0;
assign v$EXPODIFF_4412_out0 = v$MUX3_4060_out0;
assign v$ABIGGER_4745_out0 = v$ABIGGER_2412_out0;
assign v$EXPONENT_95_out0 = v$BIGGEREXPO_1814_out0;
assign v$NONVALID_424_out0 = v$NONVALID_1544_out0;
assign v$EQ8_504_out0 = v$ABSOLUTE_486_out0 == 7'h6;
assign v$EQ16_564_out0 = v$ABSOLUTE_486_out0 == 7'hc;
assign v$EQ14_785_out0 = v$ABSOLUTE_486_out0 == 7'he;
assign v$EQ13_963_out0 = v$ABSOLUTE_486_out0 == 7'hd;
assign v$EQ6_1208_out0 = v$ABSOLUTE_486_out0 == 7'h9;
assign v$EQ12_1524_out0 = v$ABSOLUTE_486_out0 == 7'h3;
assign v$G3_2173_out0 = v$ABEQUAL_341_out0 && v$Asmaller_2247_out0;
assign v$EQ7_2205_out0 = v$ABSOLUTE_486_out0 == 7'h2;
assign v$EQ9_2253_out0 = v$ABSOLUTE_486_out0 == 7'h1;
assign v$EQ2_2691_out0 = v$ABSOLUTE_486_out0 == 7'ha;
assign v$EQ1_2704_out0 = v$ABSOLUTE_486_out0 == 7'h5;
assign v$_2888_out0 = v$_1265_out1[0:0];
assign v$_2888_out1 = v$_1265_out1[9:9];
assign v$_2889_out0 = v$_1266_out1[0:0];
assign v$_2889_out1 = v$_1266_out1[9:9];
assign v$_2890_out0 = v$_1267_out1[0:0];
assign v$_2890_out1 = v$_1267_out1[9:9];
assign v$_2891_out0 = v$_1268_out1[0:0];
assign v$_2891_out1 = v$_1268_out1[9:9];
assign v$_2892_out0 = v$_1269_out1[0:0];
assign v$_2892_out1 = v$_1269_out1[9:9];
assign v$_2893_out0 = v$_1270_out1[0:0];
assign v$_2893_out1 = v$_1270_out1[9:9];
assign v$_2894_out0 = v$_1271_out1[0:0];
assign v$_2894_out1 = v$_1271_out1[9:9];
assign v$_2895_out0 = v$_1272_out1[0:0];
assign v$_2895_out1 = v$_1272_out1[9:9];
assign v$_2896_out0 = v$_1273_out1[0:0];
assign v$_2896_out1 = v$_1273_out1[9:9];
assign v$_2897_out0 = v$_1274_out1[0:0];
assign v$_2897_out1 = v$_1274_out1[9:9];
assign v$_2898_out0 = v$_1275_out1[0:0];
assign v$_2898_out1 = v$_1275_out1[9:9];
assign v$EQ5_3264_out0 = v$ABSOLUTE_486_out0 == 7'hb;
assign v$EXPODIFF_3582_out0 = v$EXPODIFF_4412_out0;
assign v$EQ11_3818_out0 = v$ABSOLUTE_486_out0 == 7'h7;
assign v$G5_3849_out0 = v$B_3507_out0 && v$_1265_out0;
assign v$G5_3850_out0 = v$B_3508_out0 && v$_1266_out0;
assign v$G5_3851_out0 = v$B_3509_out0 && v$_1267_out0;
assign v$G5_3852_out0 = v$B_3510_out0 && v$_1268_out0;
assign v$G5_3853_out0 = v$B_3511_out0 && v$_1269_out0;
assign v$G5_3854_out0 = v$B_3512_out0 && v$_1270_out0;
assign v$G5_3855_out0 = v$B_3513_out0 && v$_1271_out0;
assign v$G5_3856_out0 = v$B_3514_out0 && v$_1272_out0;
assign v$G5_3857_out0 = v$B_3515_out0 && v$_1273_out0;
assign v$G5_3858_out0 = v$B_3516_out0 && v$_1274_out0;
assign v$G5_3859_out0 = v$B_3517_out0 && v$_1275_out0;
assign v$G4_3958_out0 = v$ABEQUAL_341_out0 && v$Asmaller_2247_out0;
assign v$EQ15_4014_out0 = v$ABSOLUTE_486_out0 == 7'hf;
assign v$OP2_4043_out0 = v$OP2_2995_out0;
assign v$OP2_4044_out0 = v$OP2_2996_out0;
assign v$EQ4_4213_out0 = v$ABSOLUTE_486_out0 == 7'h0;
assign v$EQ10_5239_out0 = v$ABSOLUTE_486_out0 == 7'h8;
assign v$EQ3_5255_out0 = v$ABSOLUTE_486_out0 == 7'h4;
assign v$EXPONENT_5291_out0 = v$BIGGEREXPO_1814_out0;
assign v$10_170_out0 = v$EQ2_2691_out0;
assign v$EXPONENT_245_out0 = v$EXPODIFF_3582_out0;
assign v$3_490_out0 = v$EQ12_1524_out0;
assign v$4_718_out0 = v$EQ3_5255_out0;
assign v$13_935_out0 = v$EQ13_963_out0;
assign v$0_1011_out0 = v$EQ4_4213_out0;
assign v$MUX2_1094_out0 = v$G3_2173_out0 ? v$_3936_out0 : v$_4930_out0;
assign v$7_1310_out0 = v$EQ11_3818_out0;
assign v$6_1563_out0 = v$EQ8_504_out0;
assign v$8_1684_out0 = v$EQ10_5239_out0;
assign v$OP2_2123_out0 = v$OP2_4043_out0;
assign v$OP2_2124_out0 = v$OP2_4044_out0;
assign v$5_2475_out0 = v$EQ1_2704_out0;
assign v$_2489_out0 = v$_2888_out1[0:0];
assign v$_2489_out1 = v$_2888_out1[8:8];
assign v$_2490_out0 = v$_2889_out1[0:0];
assign v$_2490_out1 = v$_2889_out1[8:8];
assign v$_2491_out0 = v$_2890_out1[0:0];
assign v$_2491_out1 = v$_2890_out1[8:8];
assign v$_2492_out0 = v$_2891_out1[0:0];
assign v$_2492_out1 = v$_2891_out1[8:8];
assign v$_2493_out0 = v$_2892_out1[0:0];
assign v$_2493_out1 = v$_2892_out1[8:8];
assign v$_2494_out0 = v$_2893_out1[0:0];
assign v$_2494_out1 = v$_2893_out1[8:8];
assign v$_2495_out0 = v$_2894_out1[0:0];
assign v$_2495_out1 = v$_2894_out1[8:8];
assign v$_2496_out0 = v$_2895_out1[0:0];
assign v$_2496_out1 = v$_2895_out1[8:8];
assign v$_2497_out0 = v$_2896_out1[0:0];
assign v$_2497_out1 = v$_2896_out1[8:8];
assign v$_2498_out0 = v$_2897_out1[0:0];
assign v$_2498_out1 = v$_2897_out1[8:8];
assign v$_2499_out0 = v$_2898_out1[0:0];
assign v$_2499_out1 = v$_2898_out1[8:8];
assign v$12_2636_out0 = v$EQ16_564_out0;
assign v$EXPONENT_2696_out0 = v$EXPONENT_5291_out0;
assign v$G5_2945_out0 = v$G4_3958_out0 || v$ASMALLER_2055_out0;
assign v$2_3042_out0 = v$EQ7_2205_out0;
assign v$9_3255_out0 = v$EQ6_1208_out0;
assign v$MUX1_3553_out0 = v$G3_2173_out0 ? v$_4930_out0 : v$_3936_out0;
assign v$15_4218_out0 = v$EQ15_4014_out0;
assign v$14_4529_out0 = v$EQ14_785_out0;
assign v$1_4568_out0 = v$EQ9_2253_out0;
assign v$EXPONENT_4661_out0 = v$EXPONENT_95_out0;
assign v$G3_5000_out0 = v$B_3507_out0 && v$_2888_out0;
assign v$G3_5001_out0 = v$B_3508_out0 && v$_2889_out0;
assign v$G3_5002_out0 = v$B_3509_out0 && v$_2890_out0;
assign v$G3_5003_out0 = v$B_3510_out0 && v$_2891_out0;
assign v$G3_5004_out0 = v$B_3511_out0 && v$_2892_out0;
assign v$G3_5005_out0 = v$B_3512_out0 && v$_2893_out0;
assign v$G3_5006_out0 = v$B_3513_out0 && v$_2894_out0;
assign v$G3_5007_out0 = v$B_3514_out0 && v$_2895_out0;
assign v$G3_5008_out0 = v$B_3515_out0 && v$_2896_out0;
assign v$G3_5009_out0 = v$B_3516_out0 && v$_2897_out0;
assign v$G3_5010_out0 = v$B_3517_out0 && v$_2898_out0;
assign v$SEL4_275_out0 = v$EXPONENT_245_out0[3:3];
assign v$G1_373_out0 = v$12_2636_out0 || v$13_935_out0;
assign v$EQ17_719_out0 = v$EXPONENT_2696_out0 == 5'h0;
assign v$SEL3_1362_out0 = v$EXPONENT_245_out0[2:2];
assign v$XOR1_1447_out0 = v$OP2_2123_out0 ^ v$MUX1_4052_out0;
assign v$XOR1_1448_out0 = v$OP2_2124_out0 ^ v$MUX1_4053_out0;
assign v$EQ18_1971_out0 = v$EXPONENT_2696_out0 == 5'h1;
assign v$_2024_out0 = { v$EXPONENT_2696_out0,v$C19_4918_out0 };
assign v$G1_2775_out0 = v$B_3507_out0 && v$_2489_out0;
assign v$G1_2776_out0 = v$B_3508_out0 && v$_2490_out0;
assign v$G1_2777_out0 = v$B_3509_out0 && v$_2491_out0;
assign v$G1_2778_out0 = v$B_3510_out0 && v$_2492_out0;
assign v$G1_2779_out0 = v$B_3511_out0 && v$_2493_out0;
assign v$G1_2780_out0 = v$B_3512_out0 && v$_2494_out0;
assign v$G1_2781_out0 = v$B_3513_out0 && v$_2495_out0;
assign v$G1_2782_out0 = v$B_3514_out0 && v$_2496_out0;
assign v$G1_2783_out0 = v$B_3515_out0 && v$_2497_out0;
assign v$G1_2784_out0 = v$B_3516_out0 && v$_2498_out0;
assign v$G1_2785_out0 = v$B_3517_out0 && v$_2499_out0;
assign v$SMALLEREXP_3133_out0 = v$ABIGGER_4745_out0 ? v$MUX2_1094_out0 : v$MUX1_3553_out0;
assign v$LARGEREXP_3147_out0 = v$ASMALLER_2055_out0 ? v$MUX2_1094_out0 : v$MUX1_3553_out0;
assign v$_3287_out0 = { v$G5_3849_out0,v$G3_5000_out0 };
assign v$_3288_out0 = { v$G5_3850_out0,v$G3_5001_out0 };
assign v$_3289_out0 = { v$G5_3851_out0,v$G3_5002_out0 };
assign v$_3290_out0 = { v$G5_3852_out0,v$G3_5003_out0 };
assign v$_3291_out0 = { v$G5_3853_out0,v$G3_5004_out0 };
assign v$_3292_out0 = { v$G5_3854_out0,v$G3_5005_out0 };
assign v$_3293_out0 = { v$G5_3855_out0,v$G3_5006_out0 };
assign v$_3294_out0 = { v$G5_3856_out0,v$G3_5007_out0 };
assign v$_3295_out0 = { v$G5_3857_out0,v$G3_5008_out0 };
assign v$_3296_out0 = { v$G5_3858_out0,v$G3_5009_out0 };
assign v$_3297_out0 = { v$G5_3859_out0,v$G3_5010_out0 };
assign v$_3745_out0 = v$_2489_out1[0:0];
assign v$_3745_out1 = v$_2489_out1[7:7];
assign v$_3746_out0 = v$_2490_out1[0:0];
assign v$_3746_out1 = v$_2490_out1[7:7];
assign v$_3747_out0 = v$_2491_out1[0:0];
assign v$_3747_out1 = v$_2491_out1[7:7];
assign v$_3748_out0 = v$_2492_out1[0:0];
assign v$_3748_out1 = v$_2492_out1[7:7];
assign v$_3749_out0 = v$_2493_out1[0:0];
assign v$_3749_out1 = v$_2493_out1[7:7];
assign v$_3750_out0 = v$_2494_out1[0:0];
assign v$_3750_out1 = v$_2494_out1[7:7];
assign v$_3751_out0 = v$_2495_out1[0:0];
assign v$_3751_out1 = v$_2495_out1[7:7];
assign v$_3752_out0 = v$_2496_out1[0:0];
assign v$_3752_out1 = v$_2496_out1[7:7];
assign v$_3753_out0 = v$_2497_out1[0:0];
assign v$_3753_out1 = v$_2497_out1[7:7];
assign v$_3754_out0 = v$_2498_out1[0:0];
assign v$_3754_out1 = v$_2498_out1[7:7];
assign v$_3755_out0 = v$_2499_out1[0:0];
assign v$_3755_out1 = v$_2499_out1[7:7];
assign v$SWITCH_4096_out0 = v$G5_2945_out0;
assign v$B_4103_out0 = v$OP2_2123_out0;
assign v$B_4104_out0 = v$OP2_2124_out0;
assign v$G2_4494_out0 = v$14_4529_out0 || v$15_4218_out0;
assign v$SEL5_4688_out0 = v$EXPONENT_245_out0[4:4];
assign v$EQ1_4746_out0 = v$EXPONENT_4661_out0 == 5'h1e;
assign v$SEL1_4854_out0 = v$EXPONENT_245_out0[0:0];
assign v$SEL2_5204_out0 = v$EXPONENT_245_out0[1:1];
assign v$_256_out0 = v$B_4103_out0[0:0];
assign v$_256_out1 = v$B_4103_out0[15:15];
assign v$_257_out0 = v$B_4104_out0[0:0];
assign v$_257_out1 = v$B_4104_out0[15:15];
assign {v$A1_331_out1,v$A1_331_out0 } = v$OP1_1525_out0 + v$XOR1_1447_out0 + v$CIN_3082_out0;
assign {v$A1_332_out1,v$A1_332_out0 } = v$OP1_1526_out0 + v$XOR1_1448_out0 + v$CIN_3083_out0;
assign v$G16_890_out0 = v$B_3507_out0 && v$_3745_out0;
assign v$G16_891_out0 = v$B_3508_out0 && v$_3746_out0;
assign v$G16_892_out0 = v$B_3509_out0 && v$_3747_out0;
assign v$G16_893_out0 = v$B_3510_out0 && v$_3748_out0;
assign v$G16_894_out0 = v$B_3511_out0 && v$_3749_out0;
assign v$G16_895_out0 = v$B_3512_out0 && v$_3750_out0;
assign v$G16_896_out0 = v$B_3513_out0 && v$_3751_out0;
assign v$G16_897_out0 = v$B_3514_out0 && v$_3752_out0;
assign v$G16_898_out0 = v$B_3515_out0 && v$_3753_out0;
assign v$G16_899_out0 = v$B_3516_out0 && v$_3754_out0;
assign v$G16_900_out0 = v$B_3517_out0 && v$_3755_out0;
assign v$MUX4_2920_out0 = v$ABEQUAL_341_out0 ? v$MUX1_3553_out0 : v$LARGEREXP_3147_out0;
assign v$MUX22_3031_out0 = v$EQ17_719_out0 ? v$C27_3680_out0 : v$C28_1203_out0;
assign v$MUX5_3262_out0 = v$ABEQUAL_341_out0 ? v$MUX2_1094_out0 : v$SMALLEREXP_3133_out0;
assign v$G3_3467_out0 = v$G1_373_out0 || v$G2_4494_out0;
assign v$SWITCH_4809_out0 = v$SWITCH_4096_out0;
assign v$_4832_out0 = v$_3745_out1[0:0];
assign v$_4832_out1 = v$_3745_out1[6:6];
assign v$_4833_out0 = v$_3746_out1[0:0];
assign v$_4833_out1 = v$_3746_out1[6:6];
assign v$_4834_out0 = v$_3747_out1[0:0];
assign v$_4834_out1 = v$_3747_out1[6:6];
assign v$_4835_out0 = v$_3748_out1[0:0];
assign v$_4835_out1 = v$_3748_out1[6:6];
assign v$_4836_out0 = v$_3749_out1[0:0];
assign v$_4836_out1 = v$_3749_out1[6:6];
assign v$_4837_out0 = v$_3750_out1[0:0];
assign v$_4837_out1 = v$_3750_out1[6:6];
assign v$_4838_out0 = v$_3751_out1[0:0];
assign v$_4838_out1 = v$_3751_out1[6:6];
assign v$_4839_out0 = v$_3752_out1[0:0];
assign v$_4839_out1 = v$_3752_out1[6:6];
assign v$_4840_out0 = v$_3753_out1[0:0];
assign v$_4840_out1 = v$_3753_out1[6:6];
assign v$_4841_out0 = v$_3754_out1[0:0];
assign v$_4841_out1 = v$_3754_out1[6:6];
assign v$_4842_out0 = v$_3755_out1[0:0];
assign v$_4842_out1 = v$_3755_out1[6:6];
assign v$MUX23_5205_out0 = v$EQ18_1971_out0 ? v$C30_536_out0 : v$EXPONENT_2696_out0;
assign v$_11_out0 = v$_256_out1[0:0];
assign v$_11_out1 = v$_256_out1[14:14];
assign v$_12_out0 = v$_257_out1[0:0];
assign v$_12_out1 = v$_257_out1[14:14];
assign v$G1_1085_out0 = v$_4906_out0 && v$_256_out0;
assign v$G1_1086_out0 = v$_4907_out0 && v$_257_out0;
assign v$_2687_out0 = v$MUX5_3262_out0[0:0];
assign v$_2687_out1 = v$MUX5_3262_out0[11:11];
assign v$COUT_3301_out0 = v$A1_331_out1;
assign v$COUT_3302_out0 = v$A1_332_out1;
assign v$1TO4_3665_out0 = v$A1_331_out0;
assign v$1TO4_3666_out0 = v$A1_332_out0;
assign v$G4_4292_out0 = v$B_3507_out0 && v$_4832_out0;
assign v$G4_4293_out0 = v$B_3508_out0 && v$_4833_out0;
assign v$G4_4294_out0 = v$B_3509_out0 && v$_4834_out0;
assign v$G4_4295_out0 = v$B_3510_out0 && v$_4835_out0;
assign v$G4_4296_out0 = v$B_3511_out0 && v$_4836_out0;
assign v$G4_4297_out0 = v$B_3512_out0 && v$_4837_out0;
assign v$G4_4298_out0 = v$B_3513_out0 && v$_4838_out0;
assign v$G4_4299_out0 = v$B_3514_out0 && v$_4839_out0;
assign v$G4_4300_out0 = v$B_3515_out0 && v$_4840_out0;
assign v$G4_4301_out0 = v$B_3516_out0 && v$_4841_out0;
assign v$G4_4302_out0 = v$B_3517_out0 && v$_4842_out0;
assign v$_4420_out0 = v$_4832_out1[0:0];
assign v$_4420_out1 = v$_4832_out1[5:5];
assign v$_4421_out0 = v$_4833_out1[0:0];
assign v$_4421_out1 = v$_4833_out1[5:5];
assign v$_4422_out0 = v$_4834_out1[0:0];
assign v$_4422_out1 = v$_4834_out1[5:5];
assign v$_4423_out0 = v$_4835_out1[0:0];
assign v$_4423_out1 = v$_4835_out1[5:5];
assign v$_4424_out0 = v$_4836_out1[0:0];
assign v$_4424_out1 = v$_4836_out1[5:5];
assign v$_4425_out0 = v$_4837_out1[0:0];
assign v$_4425_out1 = v$_4837_out1[5:5];
assign v$_4426_out0 = v$_4838_out1[0:0];
assign v$_4426_out1 = v$_4838_out1[5:5];
assign v$_4427_out0 = v$_4839_out1[0:0];
assign v$_4427_out1 = v$_4839_out1[5:5];
assign v$_4428_out0 = v$_4840_out1[0:0];
assign v$_4428_out1 = v$_4840_out1[5:5];
assign v$_4429_out0 = v$_4841_out1[0:0];
assign v$_4429_out1 = v$_4841_out1[5:5];
assign v$_4430_out0 = v$_4842_out1[0:0];
assign v$_4430_out1 = v$_4842_out1[5:5];
assign v$G5_4434_out0 = v$SWITCH_4809_out0 && v$SUBTRACTOR_1459_out0;
assign v$G4_4572_out0 = v$EQ5_3264_out0 || v$G3_3467_out0;
assign v$_4662_out0 = { v$G1_2775_out0,v$G16_890_out0 };
assign v$_4663_out0 = { v$G1_2776_out0,v$G16_891_out0 };
assign v$_4664_out0 = { v$G1_2777_out0,v$G16_892_out0 };
assign v$_4665_out0 = { v$G1_2778_out0,v$G16_893_out0 };
assign v$_4666_out0 = { v$G1_2779_out0,v$G16_894_out0 };
assign v$_4667_out0 = { v$G1_2780_out0,v$G16_895_out0 };
assign v$_4668_out0 = { v$G1_2781_out0,v$G16_896_out0 };
assign v$_4669_out0 = { v$G1_2782_out0,v$G16_897_out0 };
assign v$_4670_out0 = { v$G1_2783_out0,v$G16_898_out0 };
assign v$_4671_out0 = { v$G1_2784_out0,v$G16_899_out0 };
assign v$_4672_out0 = { v$G1_2785_out0,v$G16_900_out0 };
assign v$_4748_out0 = v$MUX4_2920_out0[0:0];
assign v$_4748_out1 = v$MUX4_2920_out0[11:11];
assign v$G2_721_out0 = v$_1728_out0 && v$_11_out0;
assign v$G2_722_out0 = v$_1729_out0 && v$_12_out0;
assign v$TOSHIFT_1120_out0 = v$_2687_out1;
assign v$TOBIGALU_1227_out0 = v$_4748_out1;
assign v$_1940_out0 = { v$_3287_out0,v$_4662_out0 };
assign v$_1941_out0 = { v$_3288_out0,v$_4663_out0 };
assign v$_1942_out0 = { v$_3289_out0,v$_4664_out0 };
assign v$_1943_out0 = { v$_3290_out0,v$_4665_out0 };
assign v$_1944_out0 = { v$_3291_out0,v$_4666_out0 };
assign v$_1945_out0 = { v$_3292_out0,v$_4667_out0 };
assign v$_1946_out0 = { v$_3293_out0,v$_4668_out0 };
assign v$_1947_out0 = { v$_3294_out0,v$_4669_out0 };
assign v$_1948_out0 = { v$_3295_out0,v$_4670_out0 };
assign v$_1949_out0 = { v$_3296_out0,v$_4671_out0 };
assign v$_1950_out0 = { v$_3297_out0,v$_4672_out0 };
assign v$_2148_out0 = v$_4420_out1[0:0];
assign v$_2148_out1 = v$_4420_out1[4:4];
assign v$_2149_out0 = v$_4421_out1[0:0];
assign v$_2149_out1 = v$_4421_out1[4:4];
assign v$_2150_out0 = v$_4422_out1[0:0];
assign v$_2150_out1 = v$_4422_out1[4:4];
assign v$_2151_out0 = v$_4423_out1[0:0];
assign v$_2151_out1 = v$_4423_out1[4:4];
assign v$_2152_out0 = v$_4424_out1[0:0];
assign v$_2152_out1 = v$_4424_out1[4:4];
assign v$_2153_out0 = v$_4425_out1[0:0];
assign v$_2153_out1 = v$_4425_out1[4:4];
assign v$_2154_out0 = v$_4426_out1[0:0];
assign v$_2154_out1 = v$_4426_out1[4:4];
assign v$_2155_out0 = v$_4427_out1[0:0];
assign v$_2155_out1 = v$_4427_out1[4:4];
assign v$_2156_out0 = v$_4428_out1[0:0];
assign v$_2156_out1 = v$_4428_out1[4:4];
assign v$_2157_out0 = v$_4429_out1[0:0];
assign v$_2157_out1 = v$_4429_out1[4:4];
assign v$_2158_out0 = v$_4430_out1[0:0];
assign v$_2158_out1 = v$_4430_out1[4:4];
assign v$_2196_out0 = v$_11_out1[0:0];
assign v$_2196_out1 = v$_11_out1[13:13];
assign v$_2197_out0 = v$_12_out1[0:0];
assign v$_2197_out1 = v$_12_out1[13:13];
assign v$MUX8_2410_out0 = v$RET_2238_out0 ? v$C_1100_out0 : v$COUT_3301_out0;
assign v$MUX8_2411_out0 = v$RET_2239_out0 ? v$C_1101_out0 : v$COUT_3302_out0;
assign v$G15_2567_out0 = v$B_3507_out0 && v$_4420_out0;
assign v$G15_2568_out0 = v$B_3508_out0 && v$_4421_out0;
assign v$G15_2569_out0 = v$B_3509_out0 && v$_4422_out0;
assign v$G15_2570_out0 = v$B_3510_out0 && v$_4423_out0;
assign v$G15_2571_out0 = v$B_3511_out0 && v$_4424_out0;
assign v$G15_2572_out0 = v$B_3512_out0 && v$_4425_out0;
assign v$G15_2573_out0 = v$B_3513_out0 && v$_4426_out0;
assign v$G15_2574_out0 = v$B_3514_out0 && v$_4427_out0;
assign v$G15_2575_out0 = v$B_3515_out0 && v$_4428_out0;
assign v$G15_2576_out0 = v$B_3516_out0 && v$_4429_out0;
assign v$G15_2577_out0 = v$B_3517_out0 && v$_4430_out0;
assign v$SIGNTOSHIFT_3033_out0 = v$_2687_out0;
assign v$SGNBIGALU_3546_out0 = v$_4748_out0;
assign v$TOOSMALL_4217_out0 = v$G4_4572_out0;
assign v$MUX4_5267_out0 = v$G6_2973_out0 ? v$1TO4_3665_out0 : v$OP2_2123_out0;
assign v$MUX4_5268_out0 = v$G6_2974_out0 ? v$1TO4_3666_out0 : v$OP2_2124_out0;
assign v$G3_6_out0 = v$_1238_out0 && v$_2196_out0;
assign v$G3_7_out0 = v$_1239_out0 && v$_2197_out0;
assign v$SIGNTOSHIFT_255_out0 = v$SIGNTOSHIFT_3033_out0;
assign v$BIGALUSIGN_1581_out0 = v$SGNBIGALU_3546_out0;
assign v$_1701_out0 = v$_2196_out1[0:0];
assign v$_1701_out1 = v$_2196_out1[12:12];
assign v$_1702_out0 = v$_2197_out1[0:0];
assign v$_1702_out1 = v$_2197_out1[12:12];
assign v$_1912_out0 = { v$G4_4292_out0,v$G15_2567_out0 };
assign v$_1913_out0 = { v$G4_4293_out0,v$G15_2568_out0 };
assign v$_1914_out0 = { v$G4_4294_out0,v$G15_2569_out0 };
assign v$_1915_out0 = { v$G4_4295_out0,v$G15_2570_out0 };
assign v$_1916_out0 = { v$G4_4296_out0,v$G15_2571_out0 };
assign v$_1917_out0 = { v$G4_4297_out0,v$G15_2572_out0 };
assign v$_1918_out0 = { v$G4_4298_out0,v$G15_2573_out0 };
assign v$_1919_out0 = { v$G4_4299_out0,v$G15_2574_out0 };
assign v$_1920_out0 = { v$G4_4300_out0,v$G15_2575_out0 };
assign v$_1921_out0 = { v$G4_4301_out0,v$G15_2576_out0 };
assign v$_1922_out0 = { v$G4_4302_out0,v$G15_2577_out0 };
assign v$_2111_out0 = v$_2148_out1[0:0];
assign v$_2111_out1 = v$_2148_out1[3:3];
assign v$_2112_out0 = v$_2149_out1[0:0];
assign v$_2112_out1 = v$_2149_out1[3:3];
assign v$_2113_out0 = v$_2150_out1[0:0];
assign v$_2113_out1 = v$_2150_out1[3:3];
assign v$_2114_out0 = v$_2151_out1[0:0];
assign v$_2114_out1 = v$_2151_out1[3:3];
assign v$_2115_out0 = v$_2152_out1[0:0];
assign v$_2115_out1 = v$_2152_out1[3:3];
assign v$_2116_out0 = v$_2153_out1[0:0];
assign v$_2116_out1 = v$_2153_out1[3:3];
assign v$_2117_out0 = v$_2154_out1[0:0];
assign v$_2117_out1 = v$_2154_out1[3:3];
assign v$_2118_out0 = v$_2155_out1[0:0];
assign v$_2118_out1 = v$_2155_out1[3:3];
assign v$_2119_out0 = v$_2156_out1[0:0];
assign v$_2119_out1 = v$_2156_out1[3:3];
assign v$_2120_out0 = v$_2157_out1[0:0];
assign v$_2120_out1 = v$_2157_out1[3:3];
assign v$_2121_out0 = v$_2158_out1[0:0];
assign v$_2121_out1 = v$_2158_out1[3:3];
assign v$SIGNIFICANT_3533_out0 = v$TOSHIFT_1120_out0;
assign v$F1_4615_out0 = v$TOBIGALU_1227_out0;
assign v$G14_5078_out0 = v$B_3507_out0 && v$_2148_out0;
assign v$G14_5079_out0 = v$B_3508_out0 && v$_2149_out0;
assign v$G14_5080_out0 = v$B_3509_out0 && v$_2150_out0;
assign v$G14_5081_out0 = v$B_3510_out0 && v$_2151_out0;
assign v$G14_5082_out0 = v$B_3511_out0 && v$_2152_out0;
assign v$G14_5083_out0 = v$B_3512_out0 && v$_2153_out0;
assign v$G14_5084_out0 = v$B_3513_out0 && v$_2154_out0;
assign v$G14_5085_out0 = v$B_3514_out0 && v$_2155_out0;
assign v$G14_5086_out0 = v$B_3515_out0 && v$_2156_out0;
assign v$G14_5087_out0 = v$B_3516_out0 && v$_2157_out0;
assign v$G14_5088_out0 = v$B_3517_out0 && v$_2158_out0;
assign v$_5414_out0 = { v$G1_1085_out0,v$G2_721_out0 };
assign v$_5415_out0 = { v$G1_1086_out0,v$G2_722_out0 };
assign v$_350_out0 = { v$SIGNIFICANT_3533_out0,v$C12_1162_out0 };
assign v$_503_out0 = { v$SIGNIFICANT_3533_out0,v$C1_2789_out0 };
assign v$_942_out0 = { v$SIGNIFICANT_3533_out0,v$C13_1012_out0 };
assign v$_1240_out0 = { v$SIGNIFICANT_3533_out0,v$C8_598_out0 };
assign v$_1368_out0 = { v$C17_5068_out0,v$SIGNIFICANT_3533_out0 };
assign v$_1705_out0 = { v$SIGNIFICANT_3533_out0,v$C9_1514_out0 };
assign v$ASIGN_1780_out0 = v$BIGALUSIGN_1581_out0;
assign v$_2235_out0 = { v$SIGNIFICANT_3533_out0,v$C2_3117_out0 };
assign v$_2440_out0 = { v$SIGNIFICANT_3533_out0,v$C5_4307_out0 };
assign v$_2586_out0 = v$_2111_out1[0:0];
assign v$_2586_out1 = v$_2111_out1[2:2];
assign v$_2587_out0 = v$_2112_out1[0:0];
assign v$_2587_out1 = v$_2112_out1[2:2];
assign v$_2588_out0 = v$_2113_out1[0:0];
assign v$_2588_out1 = v$_2113_out1[2:2];
assign v$_2589_out0 = v$_2114_out1[0:0];
assign v$_2589_out1 = v$_2114_out1[2:2];
assign v$_2590_out0 = v$_2115_out1[0:0];
assign v$_2590_out1 = v$_2115_out1[2:2];
assign v$_2591_out0 = v$_2116_out1[0:0];
assign v$_2591_out1 = v$_2116_out1[2:2];
assign v$_2592_out0 = v$_2117_out1[0:0];
assign v$_2592_out1 = v$_2117_out1[2:2];
assign v$_2593_out0 = v$_2118_out1[0:0];
assign v$_2593_out1 = v$_2118_out1[2:2];
assign v$_2594_out0 = v$_2119_out1[0:0];
assign v$_2594_out1 = v$_2119_out1[2:2];
assign v$_2595_out0 = v$_2120_out1[0:0];
assign v$_2595_out1 = v$_2120_out1[2:2];
assign v$_2596_out0 = v$_2121_out1[0:0];
assign v$_2596_out1 = v$_2121_out1[2:2];
assign v$_2993_out0 = v$_1701_out1[0:0];
assign v$_2993_out1 = v$_1701_out1[11:11];
assign v$_2994_out0 = v$_1702_out1[0:0];
assign v$_2994_out1 = v$_1702_out1[11:11];
assign v$_3554_out0 = { v$SIGNIFICANT_3533_out0,v$C3_3005_out0 };
assign v$_3724_out0 = { v$SIGNIFICANT_3533_out0,v$C11_671_out0 };
assign v$G4_4548_out0 = v$_3126_out0 && v$_1701_out0;
assign v$G4_4549_out0 = v$_3127_out0 && v$_1702_out0;
assign v$_4579_out0 = { v$SIGNIFICANT_3533_out0,v$C7_5237_out0 };
assign v$G11_4586_out0 = v$B_3507_out0 && v$_2111_out0;
assign v$G11_4587_out0 = v$B_3508_out0 && v$_2112_out0;
assign v$G11_4588_out0 = v$B_3509_out0 && v$_2113_out0;
assign v$G11_4589_out0 = v$B_3510_out0 && v$_2114_out0;
assign v$G11_4590_out0 = v$B_3511_out0 && v$_2115_out0;
assign v$G11_4591_out0 = v$B_3512_out0 && v$_2116_out0;
assign v$G11_4592_out0 = v$B_3513_out0 && v$_2117_out0;
assign v$G11_4593_out0 = v$B_3514_out0 && v$_2118_out0;
assign v$G11_4594_out0 = v$B_3515_out0 && v$_2119_out0;
assign v$G11_4595_out0 = v$B_3516_out0 && v$_2120_out0;
assign v$G11_4596_out0 = v$B_3517_out0 && v$_2121_out0;
assign v$_4647_out0 = { v$SIGNIFICANT_3533_out0,v$C10_43_out0 };
assign v$_4683_out0 = { v$SIGNIFICANT_3533_out0,v$C4_2007_out0 };
assign v$_4752_out0 = { v$SIGNIFICANT_3533_out0,v$C6_5119_out0 };
assign v$_4828_out0 = { v$C3_4484_out0,v$F1_4615_out0 };
assign v$SIGNTOSHIFT_5047_out0 = v$SIGNTOSHIFT_255_out0;
assign v$_180_out0 = v$_2586_out1[0:0];
assign v$_180_out1 = v$_2586_out1[1:1];
assign v$_181_out0 = v$_2587_out1[0:0];
assign v$_181_out1 = v$_2587_out1[1:1];
assign v$_182_out0 = v$_2588_out1[0:0];
assign v$_182_out1 = v$_2588_out1[1:1];
assign v$_183_out0 = v$_2589_out1[0:0];
assign v$_183_out1 = v$_2589_out1[1:1];
assign v$_184_out0 = v$_2590_out1[0:0];
assign v$_184_out1 = v$_2590_out1[1:1];
assign v$_185_out0 = v$_2591_out1[0:0];
assign v$_185_out1 = v$_2591_out1[1:1];
assign v$_186_out0 = v$_2592_out1[0:0];
assign v$_186_out1 = v$_2592_out1[1:1];
assign v$_187_out0 = v$_2593_out1[0:0];
assign v$_187_out1 = v$_2593_out1[1:1];
assign v$_188_out0 = v$_2594_out1[0:0];
assign v$_188_out1 = v$_2594_out1[1:1];
assign v$_189_out0 = v$_2595_out1[0:0];
assign v$_189_out1 = v$_2595_out1[1:1];
assign v$_190_out0 = v$_2596_out1[0:0];
assign v$_190_out1 = v$_2596_out1[1:1];
assign v$2_320_out0 = v$_2235_out0;
assign v$G5_729_out0 = v$_5099_out0 && v$_2993_out0;
assign v$G5_730_out0 = v$_5100_out0 && v$_2994_out0;
assign v$_861_out0 = v$_4647_out0[8:0];
assign v$_861_out1 = v$_4647_out0[20:12];
assign v$0_1136_out0 = v$_1368_out0;
assign v$G7_1633_out0 = v$B_3507_out0 && v$_2586_out0;
assign v$G7_1634_out0 = v$B_3508_out0 && v$_2587_out0;
assign v$G7_1635_out0 = v$B_3509_out0 && v$_2588_out0;
assign v$G7_1636_out0 = v$B_3510_out0 && v$_2589_out0;
assign v$G7_1637_out0 = v$B_3511_out0 && v$_2590_out0;
assign v$G7_1638_out0 = v$B_3512_out0 && v$_2591_out0;
assign v$G7_1639_out0 = v$B_3513_out0 && v$_2592_out0;
assign v$G7_1640_out0 = v$B_3514_out0 && v$_2593_out0;
assign v$G7_1641_out0 = v$B_3515_out0 && v$_2594_out0;
assign v$G7_1642_out0 = v$B_3516_out0 && v$_2595_out0;
assign v$G7_1643_out0 = v$B_3517_out0 && v$_2596_out0;
assign v$_1812_out0 = v$_4579_out0[5:0];
assign v$_1812_out1 = v$_4579_out0[17:12];
assign v$_1871_out0 = v$_4752_out0[4:0];
assign v$_1871_out1 = v$_4752_out0[16:12];
assign v$_2401_out0 = v$_350_out0[10:0];
assign v$_2401_out1 = v$_350_out0[22:12];
assign v$_2428_out0 = v$_4683_out0[2:0];
assign v$_2428_out1 = v$_4683_out0[14:12];
assign v$_2639_out0 = v$_1240_out0[6:0];
assign v$_2639_out1 = v$_1240_out0[18:12];
assign v$_2750_out0 = { v$C15_3806_out0,v$_503_out0 };
assign v$_3125_out0 = v$_1705_out0[7:0];
assign v$_3125_out1 = v$_1705_out0[19:12];
assign v$_3221_out0 = { v$G14_5078_out0,v$G11_4586_out0 };
assign v$_3222_out0 = { v$G14_5079_out0,v$G11_4587_out0 };
assign v$_3223_out0 = { v$G14_5080_out0,v$G11_4588_out0 };
assign v$_3224_out0 = { v$G14_5081_out0,v$G11_4589_out0 };
assign v$_3225_out0 = { v$G14_5082_out0,v$G11_4590_out0 };
assign v$_3226_out0 = { v$G14_5083_out0,v$G11_4591_out0 };
assign v$_3227_out0 = { v$G14_5084_out0,v$G11_4592_out0 };
assign v$_3228_out0 = { v$G14_5085_out0,v$G11_4593_out0 };
assign v$_3229_out0 = { v$G14_5086_out0,v$G11_4594_out0 };
assign v$_3230_out0 = { v$G14_5087_out0,v$G11_4595_out0 };
assign v$_3231_out0 = { v$G14_5088_out0,v$G11_4596_out0 };
assign v$_3366_out0 = v$_3554_out0[1:0];
assign v$_3366_out1 = v$_3554_out0[13:12];
assign v$_3549_out0 = v$_942_out0[11:0];
assign v$_3549_out1 = v$_942_out0[23:12];
assign v$G6_3552_out0 = ! v$ASIGN_1780_out0;
assign v$_3807_out0 = v$_3724_out0[9:0];
assign v$_3807_out1 = v$_3724_out0[21:12];
assign v$_3877_out0 = { v$G3_6_out0,v$G4_4548_out0 };
assign v$_3878_out0 = { v$G3_7_out0,v$G4_4549_out0 };
assign v$_4820_out0 = v$_2993_out1[0:0];
assign v$_4820_out1 = v$_2993_out1[10:10];
assign v$_4821_out0 = v$_2994_out1[0:0];
assign v$_4821_out1 = v$_2994_out1[10:10];
assign v$_4870_out0 = v$_2440_out0[3:0];
assign v$_4870_out1 = v$_2440_out0[15:12];
assign v$MUX3_693_out0 = v$G5_4434_out0 ? v$G6_3552_out0 : v$ASIGN_1780_out0;
assign v$EQ9_901_out0 = v$_3807_out0 == 10'h0;
assign v$EQ11_1119_out0 = v$_3549_out0 == 12'h0;
assign v$1_2087_out0 = v$_2750_out0;
assign v$G12_2209_out0 = v$B_3507_out0 && v$_180_out0;
assign v$G12_2210_out0 = v$B_3508_out0 && v$_181_out0;
assign v$G12_2211_out0 = v$B_3509_out0 && v$_182_out0;
assign v$G12_2212_out0 = v$B_3510_out0 && v$_183_out0;
assign v$G12_2213_out0 = v$B_3511_out0 && v$_184_out0;
assign v$G12_2214_out0 = v$B_3512_out0 && v$_185_out0;
assign v$G12_2215_out0 = v$B_3513_out0 && v$_186_out0;
assign v$G12_2216_out0 = v$B_3514_out0 && v$_187_out0;
assign v$G12_2217_out0 = v$B_3515_out0 && v$_188_out0;
assign v$G12_2218_out0 = v$B_3516_out0 && v$_189_out0;
assign v$G12_2219_out0 = v$B_3517_out0 && v$_190_out0;
assign v$_2342_out0 = { v$_1912_out0,v$_3221_out0 };
assign v$_2343_out0 = { v$_1913_out0,v$_3222_out0 };
assign v$_2344_out0 = { v$_1914_out0,v$_3223_out0 };
assign v$_2345_out0 = { v$_1915_out0,v$_3224_out0 };
assign v$_2346_out0 = { v$_1916_out0,v$_3225_out0 };
assign v$_2347_out0 = { v$_1917_out0,v$_3226_out0 };
assign v$_2348_out0 = { v$_1918_out0,v$_3227_out0 };
assign v$_2349_out0 = { v$_1919_out0,v$_3228_out0 };
assign v$_2350_out0 = { v$_1920_out0,v$_3229_out0 };
assign v$_2351_out0 = { v$_1921_out0,v$_3230_out0 };
assign v$_2352_out0 = { v$_1922_out0,v$_3231_out0 };
assign v$_2620_out0 = { v$_5414_out0,v$_3877_out0 };
assign v$_2621_out0 = { v$_5415_out0,v$_3878_out0 };
assign v$_2670_out0 = v$_4820_out1[0:0];
assign v$_2670_out1 = v$_4820_out1[9:9];
assign v$_2671_out0 = v$_4821_out1[0:0];
assign v$_2671_out1 = v$_4821_out1[9:9];
assign v$EQ7_2953_out0 = v$_3125_out0 == 8'h0;
assign v$EQ2_3106_out0 = v$_2428_out0 == 3'h0;
assign v$G6_3165_out0 = v$B_3507_out0 && v$_180_out1;
assign v$G6_3166_out0 = v$B_3508_out0 && v$_181_out1;
assign v$G6_3167_out0 = v$B_3509_out0 && v$_182_out1;
assign v$G6_3168_out0 = v$B_3510_out0 && v$_183_out1;
assign v$G6_3169_out0 = v$B_3511_out0 && v$_184_out1;
assign v$G6_3170_out0 = v$B_3512_out0 && v$_185_out1;
assign v$G6_3171_out0 = v$B_3513_out0 && v$_186_out1;
assign v$G6_3172_out0 = v$B_3514_out0 && v$_187_out1;
assign v$G6_3173_out0 = v$B_3515_out0 && v$_188_out1;
assign v$G6_3174_out0 = v$B_3516_out0 && v$_189_out1;
assign v$G6_3175_out0 = v$B_3517_out0 && v$_190_out1;
assign v$EQ1_3286_out0 = v$_3366_out0 == 2'h0;
assign v$EQ8_3440_out0 = v$_861_out0 == 9'h0;
assign v$EQ3_3655_out0 = v$_4870_out0 == 4'h0;
assign v$EQ5_3791_out0 = v$_1812_out0 == 6'h0;
assign v$EQ10_3887_out0 = v$_2401_out0 == 11'h0;
assign v$G6_4354_out0 = v$_4723_out0 && v$_4820_out0;
assign v$G6_4355_out0 = v$_4724_out0 && v$_4821_out0;
assign v$EQ6_4783_out0 = v$_2639_out0 == 7'h0;
assign v$EQ4_5183_out0 = v$_1871_out0 == 5'h0;
assign v$G10_59_out0 = ! v$EQ10_3887_out0;
assign v$G9_91_out0 = ! v$EQ9_901_out0;
assign v$_118_out0 = { v$G7_1633_out0,v$G12_2209_out0 };
assign v$_119_out0 = { v$G7_1634_out0,v$G12_2210_out0 };
assign v$_120_out0 = { v$G7_1635_out0,v$G12_2211_out0 };
assign v$_121_out0 = { v$G7_1636_out0,v$G12_2212_out0 };
assign v$_122_out0 = { v$G7_1637_out0,v$G12_2213_out0 };
assign v$_123_out0 = { v$G7_1638_out0,v$G12_2214_out0 };
assign v$_124_out0 = { v$G7_1639_out0,v$G12_2215_out0 };
assign v$_125_out0 = { v$G7_1640_out0,v$G12_2216_out0 };
assign v$_126_out0 = { v$G7_1641_out0,v$G12_2217_out0 };
assign v$_127_out0 = { v$G7_1642_out0,v$G12_2218_out0 };
assign v$_128_out0 = { v$G7_1643_out0,v$G12_2219_out0 };
assign v$G4_1102_out0 = ! v$EQ4_5183_out0;
assign v$G2_1233_out0 = ! v$EQ2_3106_out0;
assign v$_1644_out0 = { v$_1940_out0,v$_2342_out0 };
assign v$_1645_out0 = { v$_1941_out0,v$_2343_out0 };
assign v$_1646_out0 = { v$_1942_out0,v$_2344_out0 };
assign v$_1647_out0 = { v$_1943_out0,v$_2345_out0 };
assign v$_1648_out0 = { v$_1944_out0,v$_2346_out0 };
assign v$_1649_out0 = { v$_1945_out0,v$_2347_out0 };
assign v$_1650_out0 = { v$_1946_out0,v$_2348_out0 };
assign v$_1651_out0 = { v$_1947_out0,v$_2349_out0 };
assign v$_1652_out0 = { v$_1948_out0,v$_2350_out0 };
assign v$_1653_out0 = { v$_1949_out0,v$_2351_out0 };
assign v$_1654_out0 = { v$_1950_out0,v$_2352_out0 };
assign v$G6_2012_out0 = ! v$EQ6_4783_out0;
assign v$G8_2419_out0 = ! v$EQ8_3440_out0;
assign v$_2711_out0 = { v$G5_729_out0,v$G6_4354_out0 };
assign v$_2712_out0 = { v$G5_730_out0,v$G6_4355_out0 };
assign v$G7_2835_out0 = ! v$EQ7_2953_out0;
assign v$G1_3684_out0 = ! v$EQ1_3286_out0;
assign v$MUX1_3727_out0 = v$SEL1_4854_out0 ? v$1_2087_out0 : v$0_1136_out0;
assign v$G7_3779_out0 = v$_5048_out0 && v$_2670_out0;
assign v$G7_3780_out0 = v$_5049_out0 && v$_2671_out0;
assign v$G5_4111_out0 = ! v$EQ5_3791_out0;
assign v$_4349_out0 = v$_2670_out1[0:0];
assign v$_4349_out1 = v$_2670_out1[8:8];
assign v$_4350_out0 = v$_2671_out1[0:0];
assign v$_4350_out1 = v$_2671_out1[8:8];
assign v$SIGN_5044_out0 = v$MUX3_693_out0;
assign v$G11_5397_out0 = ! v$EQ11_1119_out0;
assign v$G3_5425_out0 = ! v$EQ3_3655_out0;
assign v$_164_out0 = { v$G10_59_out0,v$_2401_out1 };
assign v$_607_out0 = { v$G6_2012_out0,v$_2639_out1 };
assign v$NOTUSE12_947_out0 = v$G10_59_out0;
assign v$SIGN_1005_out0 = v$SIGN_5044_out0;
assign v$_1523_out0 = { v$G7_2835_out0,v$_3125_out1 };
assign v$_1549_out0 = { v$G4_1102_out0,v$_1871_out1 };
assign v$NOTUSE4_1839_out0 = v$G2_1233_out0;
assign v$_2027_out0 = { v$G2_1233_out0,v$_2428_out1 };
assign v$NOTUSE10_2286_out0 = v$G8_2419_out0;
assign v$NOTUSE7_2361_out0 = v$G5_4111_out0;
assign v$_2501_out0 = { v$G9_91_out0,v$_3807_out1 };
assign v$_2637_out0 = { v$G5_4111_out0,v$_1812_out1 };
assign v$NOTUSE6_2721_out0 = v$G4_1102_out0;
assign v$_2760_out0 = v$_4349_out1[0:0];
assign v$_2760_out1 = v$_4349_out1[7:7];
assign v$_2761_out0 = v$_4350_out1[0:0];
assign v$_2761_out1 = v$_4350_out1[7:7];
assign v$G8_2899_out0 = v$_2378_out0 && v$_4349_out0;
assign v$G8_2900_out0 = v$_2379_out0 && v$_4350_out0;
assign v$_3000_out0 = { v$G3_5425_out0,v$_4870_out1 };
assign v$_3050_out0 = { v$G11_5397_out0,v$_3549_out1 };
assign v$NOTUSE13_3468_out0 = v$G11_5397_out0;
assign v$NOTUSE11_3709_out0 = v$G9_91_out0;
assign v$_3860_out0 = { v$G1_3684_out0,v$_3366_out1 };
assign v$_3901_out0 = { v$G8_2419_out0,v$_861_out1 };
assign v$NOTUSE5_3950_out0 = v$G3_5425_out0;
assign v$NOTUSE8_5140_out0 = v$G6_2012_out0;
assign v$NOTUSE9_5190_out0 = v$G7_2835_out0;
assign v$_5433_out0 = { v$_118_out0,v$G6_3165_out0 };
assign v$_5434_out0 = { v$_119_out0,v$G6_3166_out0 };
assign v$_5435_out0 = { v$_120_out0,v$G6_3167_out0 };
assign v$_5436_out0 = { v$_121_out0,v$G6_3168_out0 };
assign v$_5437_out0 = { v$_122_out0,v$G6_3169_out0 };
assign v$_5438_out0 = { v$_123_out0,v$G6_3170_out0 };
assign v$_5439_out0 = { v$_124_out0,v$G6_3171_out0 };
assign v$_5440_out0 = { v$_125_out0,v$G6_3172_out0 };
assign v$_5441_out0 = { v$_126_out0,v$G6_3173_out0 };
assign v$_5442_out0 = { v$_127_out0,v$G6_3174_out0 };
assign v$_5443_out0 = { v$_128_out0,v$G6_3175_out0 };
assign v$7_129_out0 = v$_2637_out0;
assign v$13_273_out0 = v$_3050_out0;
assign v$5_428_out0 = v$_3000_out0;
assign v$12_499_out0 = v$_164_out0;
assign v$4_989_out0 = v$_2027_out0;
assign v$_1188_out0 = { v$_1644_out0,v$_5433_out0 };
assign v$_1189_out0 = { v$_1645_out0,v$_5434_out0 };
assign v$_1190_out0 = { v$_1646_out0,v$_5435_out0 };
assign v$_1191_out0 = { v$_1647_out0,v$_5436_out0 };
assign v$_1192_out0 = { v$_1648_out0,v$_5437_out0 };
assign v$_1193_out0 = { v$_1649_out0,v$_5438_out0 };
assign v$_1194_out0 = { v$_1650_out0,v$_5439_out0 };
assign v$_1195_out0 = { v$_1651_out0,v$_5440_out0 };
assign v$_1196_out0 = { v$_1652_out0,v$_5441_out0 };
assign v$_1197_out0 = { v$_1653_out0,v$_5442_out0 };
assign v$_1198_out0 = { v$_1654_out0,v$_5443_out0 };
assign v$3_1416_out0 = v$_3860_out0;
assign v$G9_1426_out0 = v$_4250_out0 && v$_2760_out0;
assign v$G9_1427_out0 = v$_4251_out0 && v$_2761_out0;
assign v$_1720_out0 = { v$G7_3779_out0,v$G8_2899_out0 };
assign v$_1721_out0 = { v$G7_3780_out0,v$G8_2900_out0 };
assign v$NEWSIGN_3096_out0 = v$SIGN_1005_out0;
assign v$9_3469_out0 = v$_1523_out0;
assign v$6_3566_out0 = v$_1549_out0;
assign v$11_3593_out0 = v$_2501_out0;
assign v$8_3965_out0 = v$_607_out0;
assign v$_4633_out0 = v$_2760_out1[0:0];
assign v$_4633_out1 = v$_2760_out1[6:6];
assign v$_4634_out0 = v$_2761_out1[0:0];
assign v$_4634_out1 = v$_2761_out1[6:6];
assign v$10_4736_out0 = v$_3901_out0;
assign v$_242_out0 = v$_4633_out1[0:0];
assign v$_242_out1 = v$_4633_out1[5:5];
assign v$_243_out0 = v$_4634_out1[0:0];
assign v$_243_out1 = v$_4634_out1[5:5];
assign v$X1_381_out0 = v$_1188_out0;
assign v$X1_382_out0 = v$_1189_out0;
assign v$X1_383_out0 = v$_1190_out0;
assign v$X1_384_out0 = v$_1191_out0;
assign v$X1_385_out0 = v$_1192_out0;
assign v$X1_386_out0 = v$_1193_out0;
assign v$X1_387_out0 = v$_1194_out0;
assign v$X1_388_out0 = v$_1195_out0;
assign v$X1_389_out0 = v$_1196_out0;
assign v$X1_390_out0 = v$_1197_out0;
assign v$X1_391_out0 = v$_1198_out0;
assign v$_399_out0 = { v$_2711_out0,v$_1720_out0 };
assign v$_400_out0 = { v$_2712_out0,v$_1721_out0 };
assign v$G10_2910_out0 = v$_2717_out0 && v$_4633_out0;
assign v$G10_2911_out0 = v$_2718_out0 && v$_4634_out0;
assign v$MUX3_3189_out0 = v$SEL1_4854_out0 ? v$5_428_out0 : v$4_989_out0;
assign v$MUX5_3232_out0 = v$SEL1_4854_out0 ? v$9_3469_out0 : v$8_3965_out0;
assign v$MUX4_3470_out0 = v$SEL1_4854_out0 ? v$7_129_out0 : v$6_3566_out0;
assign v$MUX7_3999_out0 = v$SEL1_4854_out0 ? v$13_273_out0 : v$12_499_out0;
assign v$MUX2_4855_out0 = v$SEL1_4854_out0 ? v$3_1416_out0 : v$2_320_out0;
assign v$MUX6_5236_out0 = v$SEL1_4854_out0 ? v$11_3593_out0 : v$10_4736_out0;
assign v$_8_out0 = { v$C8_4137_out0,v$X1_390_out0 };
assign v$B0_90_out0 = v$X1_382_out0;
assign v$_104_out0 = { v$C10_2703_out0,v$X1_381_out0 };
assign v$_517_out0 = { v$C5_1899_out0,v$X1_389_out0 };
assign v$_708_out0 = { v$C9_3863_out0,v$X1_388_out0 };
assign v$_745_out0 = { v$_2620_out0,v$_399_out0 };
assign v$_746_out0 = { v$_2621_out0,v$_400_out0 };
assign v$_950_out0 = { v$C7_4637_out0,v$X1_386_out0 };
assign v$MUX14_1305_out0 = v$SEL2_5204_out0 ? v$C18_2405_out0 : v$MUX7_3999_out0;
assign v$G11_1316_out0 = v$_5027_out0 && v$_242_out0;
assign v$G11_1317_out0 = v$_5028_out0 && v$_243_out0;
assign v$_1411_out0 = { v$C2_2749_out0,v$X1_384_out0 };
assign v$_1449_out0 = { v$C4_777_out0,v$X1_391_out0 };
assign v$MUX10_1481_out0 = v$SEL2_5204_out0 ? v$MUX6_5236_out0 : v$MUX5_3232_out0;
assign v$_2069_out0 = { v$C1_3612_out0,v$X1_383_out0 };
assign v$MUX8_2088_out0 = v$SEL2_5204_out0 ? v$MUX2_4855_out0 : v$MUX1_3727_out0;
assign v$_2623_out0 = v$_242_out1[0:0];
assign v$_2623_out1 = v$_242_out1[4:4];
assign v$_2624_out0 = v$_243_out1[0:0];
assign v$_2624_out1 = v$_243_out1[4:4];
assign v$_3792_out0 = { v$C3_4571_out0,v$X1_387_out0 };
assign v$_4270_out0 = { v$G9_1426_out0,v$G10_2910_out0 };
assign v$_4271_out0 = { v$G9_1427_out0,v$G10_2911_out0 };
assign v$MUX9_4512_out0 = v$SEL2_5204_out0 ? v$MUX4_3470_out0 : v$MUX3_3189_out0;
assign v$_5390_out0 = { v$C6_3524_out0,v$X1_385_out0 };
assign v$B6_262_out0 = v$_5390_out0;
assign v$B10_317_out0 = v$_708_out0;
assign v$B4_380_out0 = v$_517_out0;
assign v$B3_692_out0 = v$_3792_out0;
assign v$B7_1140_out0 = v$_104_out0;
assign v$B2_1666_out0 = v$_1411_out0;
assign v$B9_1681_out0 = v$_950_out0;
assign v$B8_2200_out0 = v$_8_out0;
assign v$B1_2488_out0 = v$_2069_out0;
assign v$B5_2508_out0 = v$_1449_out0;
assign v$MUX11_2798_out0 = v$SEL3_1362_out0 ? v$MUX9_4512_out0 : v$MUX8_2088_out0;
assign v$_2949_out0 = v$_2623_out1[0:0];
assign v$_2949_out1 = v$_2623_out1[3:3];
assign v$_2950_out0 = v$_2624_out1[0:0];
assign v$_2950_out1 = v$_2624_out1[3:3];
assign v$G12_3199_out0 = v$_1297_out0 && v$_2623_out0;
assign v$G12_3200_out0 = v$_1298_out0 && v$_2624_out0;
assign v$MUX12_3802_out0 = v$SEL3_1362_out0 ? v$MUX14_1305_out0 : v$MUX10_1481_out0;
assign v$B0_4321_out0 = v$B0_90_out0;
assign v$_773_out0 = v$_2949_out1[0:0];
assign v$_773_out1 = v$_2949_out1[2:2];
assign v$_774_out0 = v$_2950_out1[0:0];
assign v$_774_out1 = v$_2950_out1[2:2];
assign v$B9_812_out0 = v$B9_1681_out0;
assign v$B2_1401_out0 = v$B2_1666_out0;
assign v$SEL3_1892_out0 = v$B0_4321_out0[1:1];
assign v$B8_1901_out0 = v$B8_2200_out0;
assign v$G13_2037_out0 = v$_4804_out0 && v$_2949_out0;
assign v$G13_2038_out0 = v$_4805_out0 && v$_2950_out0;
assign v$B6_2056_out0 = v$B6_262_out0;
assign v$B7_3060_out0 = v$B7_1140_out0;
assign v$B5_3091_out0 = v$B5_2508_out0;
assign v$B3_3095_out0 = v$B3_692_out0;
assign v$MUX13_3550_out0 = v$SEL4_275_out0 ? v$MUX12_3802_out0 : v$MUX11_2798_out0;
assign v$SEL16_3804_out0 = v$B0_4321_out0[10:2];
assign v$B4_4037_out0 = v$B4_380_out0;
assign v$B10_4097_out0 = v$B10_317_out0;
assign v$B1_4597_out0 = v$B1_2488_out0;
assign v$SEL1_4808_out0 = v$B0_4321_out0[0:0];
assign v$_4968_out0 = { v$G11_1316_out0,v$G12_3199_out0 };
assign v$_4969_out0 = { v$G11_1317_out0,v$G12_3200_out0 };
assign v$SEL28_143_out0 = v$B4_4037_out0[4:4];
assign v$G14_285_out0 = v$_223_out0 && v$_773_out0;
assign v$G14_286_out0 = v$_224_out0 && v$_774_out0;
assign v$SEL22_514_out0 = v$B4_4037_out0[14:14];
assign v$SEL26_529_out0 = v$B5_3091_out0[15:15];
assign v$SEL32_696_out0 = v$B7_3060_out0[17:17];
assign v$SEL39_727_out0 = v$B8_1901_out0[16:8];
assign v$SEL20_848_out0 = v$B1_4597_out0[11:11];
assign v$SEL37_997_out0 = v$B7_3060_out0[16:8];
assign v$SEL18_1412_out0 = v$B2_1401_out0[10:2];
assign v$SEL35_1547_out0 = v$B6_2056_out0[6:6];
assign v$SEL33_1822_out0 = v$B8_1901_out0[18:18];
assign v$SEL17_1907_out0 = v$B1_4597_out0[10:2];
assign v$SEL24_2372_out0 = v$B3_3095_out0[4:4];
assign v$SEL36_2407_out0 = v$B6_2056_out0[16:8];
assign v$SEL34_2547_out0 = v$B6_2056_out0[7:7];
assign v$SEL30_2716_out0 = v$B3_3095_out0[3:3];
assign v$SEL27_2724_out0 = v$B3_3095_out0[13:5];
assign v$SEL21_2848_out0 = v$B2_1401_out0[12:12];
assign v$SEL86_2965_out0 = v$B10_4097_out0[19:10];
assign v$SEL25_3032_out0 = v$B4_4037_out0[13:5];
assign v$SEL85_3247_out0 = v$B9_812_out0[19:10];
assign v$_3591_out0 = { v$_4270_out0,v$_4968_out0 };
assign v$_3592_out0 = { v$_4271_out0,v$_4969_out0 };
assign v$C_3603_out0 = v$SEL16_3804_out0;
assign v$SEL84_4290_out0 = v$B9_812_out0[9:9];
assign v$SEL2_4366_out0 = v$B1_4597_out0[1:1];
assign v$SEL29_4456_out0 = v$B5_3091_out0[14:14];
assign v$SEL38_4463_out0 = v$B8_1901_out0[17:17];
assign v$SEL88_4558_out0 = v$B10_4097_out0[20:20];
assign v$SEL31_4563_out0 = v$B7_3060_out0[7:7];
assign v$SEL23_4774_out0 = v$B5_3091_out0[13:5];
assign v$SEL19_4778_out0 = v$B2_1401_out0[11:11];
assign v$A_4976_out0 = v$SEL3_1892_out0;
assign v$_5143_out0 = v$_773_out1[0:0];
assign v$_5143_out1 = v$_773_out1[1:1];
assign v$_5144_out0 = v$_774_out1[0:0];
assign v$_5144_out1 = v$_774_out1[1:1];
assign v$MUX15_5166_out0 = v$SEL5_4688_out0 ? v$C18_2405_out0 : v$MUX13_3550_out0;
assign v$B_61_out0 = v$SEL28_143_out0;
assign v$B_63_out0 = v$SEL84_4290_out0;
assign v$B_66_out0 = v$SEL2_4366_out0;
assign v$B_67_out0 = v$SEL22_514_out0;
assign v$B_72_out0 = v$SEL20_848_out0;
assign v$B_73_out0 = v$SEL32_696_out0;
assign v$B_77_out0 = v$SEL31_4563_out0;
assign v$_272_out0 = { v$C3_4882_out0,v$SEL30_2716_out0 };
assign v$SEL21_756_out0 = v$C_3603_out0[1:1];
assign v$SEL22_960_out0 = v$C_3603_out0[5:5];
assign v$SEL19_1488_out0 = v$C_3603_out0[4:4];
assign v$SEL26_1708_out0 = v$C_3603_out0[8:8];
assign v$SEL24_1793_out0 = v$C_3603_out0[3:3];
assign v$G16_1803_out0 = v$_1512_out1 && v$_5143_out1;
assign v$G16_1804_out0 = v$_1513_out1 && v$_5144_out1;
assign v$G15_2300_out0 = v$_1512_out0 && v$_5143_out0;
assign v$G15_2301_out0 = v$_1513_out0 && v$_5144_out0;
assign v$SEL27_2609_out0 = v$C_3603_out0[7:7];
assign v$G3_2808_out0 = ! v$A_4976_out0;
assign v$_3547_out0 = { v$G13_2037_out0,v$G14_285_out0 };
assign v$_3548_out0 = { v$G13_2038_out0,v$G14_286_out0 };
assign v$A_3570_out0 = v$SEL85_3247_out0;
assign v$C_3602_out0 = v$SEL27_2724_out0;
assign v$C_3604_out0 = v$SEL36_2407_out0;
assign v$A_3705_out0 = v$SEL23_4774_out0;
assign v$A_3706_out0 = v$SEL18_1412_out0;
assign v$A_3707_out0 = v$SEL39_727_out0;
assign v$B_3712_out0 = v$SEL25_3032_out0;
assign v$B_3713_out0 = v$SEL17_1907_out0;
assign v$B_3714_out0 = v$SEL37_997_out0;
assign v$SEL23_3970_out0 = v$C_3603_out0[6:6];
assign v$C_4519_out0 = v$SEL86_2965_out0;
assign v$SEL20_4545_out0 = v$C_3603_out0[0:0];
assign v$SEL25_4657_out0 = v$C_3603_out0[2:2];
assign v$A_4971_out0 = v$SEL24_2372_out0;
assign v$A_4977_out0 = v$SEL29_4456_out0;
assign v$A_4982_out0 = v$SEL19_4778_out0;
assign v$A_4983_out0 = v$SEL38_4463_out0;
assign v$A_4987_out0 = v$SEL34_2547_out0;
assign v$SHIFTSIGNIFICANT_5041_out0 = v$MUX15_5166_out0;
assign v$_5429_out0 = { v$C5_2191_out0,v$SEL35_1547_out0 };
assign v$SEL4_40_out0 = v$C_4519_out0[5:5];
assign v$SEL3_358_out0 = v$A_3705_out0[4:4];
assign v$SEL3_359_out0 = v$A_3706_out0[4:4];
assign v$SEL3_360_out0 = v$A_3707_out0[4:4];
assign v$SEL2_605_out0 = v$A_3570_out0[6:6];
assign v$SEL2_740_out0 = v$A_3705_out0[6:6];
assign v$SEL2_741_out0 = v$A_3706_out0[6:6];
assign v$SEL2_742_out0 = v$A_3707_out0[6:6];
assign v$SEL21_755_out0 = v$C_3602_out0[1:1];
assign v$SEL21_757_out0 = v$C_3604_out0[1:1];
assign v$SEL15_832_out0 = v$A_3570_out0[2:2];
assign v$SEL27_919_out0 = v$A_3570_out0[3:3];
assign v$SEL22_959_out0 = v$C_3602_out0[5:5];
assign v$SEL22_961_out0 = v$C_3604_out0[5:5];
assign v$SEL17_994_out0 = v$A_3570_out0[0:0];
assign v$SEL6_1042_out0 = v$A_3705_out0[5:5];
assign v$SEL6_1043_out0 = v$A_3706_out0[5:5];
assign v$SEL6_1044_out0 = v$A_3707_out0[5:5];
assign v$SEL10_1159_out0 = v$B_3712_out0[4:4];
assign v$SEL10_1160_out0 = v$B_3713_out0[4:4];
assign v$SEL10_1161_out0 = v$B_3714_out0[4:4];
assign v$G4_1331_out0 = ! v$B_61_out0;
assign v$G4_1333_out0 = ! v$B_63_out0;
assign v$G4_1336_out0 = ! v$B_66_out0;
assign v$G4_1337_out0 = ! v$B_67_out0;
assign v$G4_1342_out0 = ! v$B_72_out0;
assign v$G4_1343_out0 = ! v$B_73_out0;
assign v$G4_1347_out0 = ! v$B_77_out0;
assign v$SEL15_1364_out0 = v$B_3712_out0[0:0];
assign v$SEL15_1365_out0 = v$B_3713_out0[0:0];
assign v$SEL15_1366_out0 = v$B_3714_out0[0:0];
assign v$SEL24_1409_out0 = v$C_4519_out0[0:0];
assign v$SEL19_1487_out0 = v$C_3602_out0[4:4];
assign v$SEL19_1489_out0 = v$C_3604_out0[4:4];
assign v$SEL14_1492_out0 = v$B_3712_out0[1:1];
assign v$SEL14_1493_out0 = v$B_3713_out0[1:1];
assign v$SEL14_1494_out0 = v$B_3714_out0[1:1];
assign v$SEL8_1505_out0 = v$C_4519_out0[4:4];
assign v$SEL30_1615_out0 = v$C_4519_out0[9:9];
assign v$SEL3_1664_out0 = v$C_4519_out0[1:1];
assign v$SEL26_1707_out0 = v$C_3602_out0[8:8];
assign v$SEL26_1709_out0 = v$C_3604_out0[8:8];
assign v$SEL26_1765_out0 = v$A_3570_out0[7:7];
assign v$SEL24_1792_out0 = v$C_3602_out0[3:3];
assign v$SEL24_1794_out0 = v$C_3604_out0[3:3];
assign v$SEL16_1897_out0 = v$A_3570_out0[1:1];
assign v$SEL12_2082_out0 = v$B_3712_out0[5:5];
assign v$SEL12_2083_out0 = v$B_3713_out0[5:5];
assign v$SEL12_2084_out0 = v$B_3714_out0[5:5];
assign v$C7_2319_out0 = v$SEL27_2609_out0;
assign v$G1_2523_out0 = v$G3_2808_out0 && v$B_66_out0;
assign v$SEL11_2550_out0 = v$B_3712_out0[6:6];
assign v$SEL11_2551_out0 = v$B_3713_out0[6:6];
assign v$SEL11_2552_out0 = v$B_3714_out0[6:6];
assign v$SEL27_2608_out0 = v$C_3602_out0[7:7];
assign v$SEL27_2610_out0 = v$C_3604_out0[7:7];
assign v$C6_2676_out0 = v$SEL23_3970_out0;
assign v$G3_2803_out0 = ! v$A_4971_out0;
assign v$G3_2809_out0 = ! v$A_4977_out0;
assign v$G3_2814_out0 = ! v$A_4982_out0;
assign v$G3_2815_out0 = ! v$A_4983_out0;
assign v$G3_2819_out0 = ! v$A_4987_out0;
assign v$SEL22_2924_out0 = v$A_3570_out0[8:8];
assign v$SEL11_3136_out0 = v$C_4519_out0[3:3];
assign v$SEL4_3162_out0 = v$A_3705_out0[2:2];
assign v$SEL4_3163_out0 = v$A_3706_out0[2:2];
assign v$SEL4_3164_out0 = v$A_3707_out0[2:2];
assign v$SEL1_3203_out0 = v$A_3570_out0[4:4];
assign v$SEL1_3306_out0 = v$A_3705_out0[1:1];
assign v$SEL1_3307_out0 = v$A_3706_out0[1:1];
assign v$SEL1_3308_out0 = v$A_3707_out0[1:1];
assign v$SEL9_3387_out0 = v$A_3705_out0[0:0];
assign v$SEL9_3388_out0 = v$A_3706_out0[0:0];
assign v$SEL9_3389_out0 = v$A_3707_out0[0:0];
assign v$C4_3420_out0 = v$SEL19_1488_out0;
assign v$SEL18_3450_out0 = v$B_3712_out0[3:3];
assign v$SEL18_3451_out0 = v$B_3713_out0[3:3];
assign v$SEL18_3452_out0 = v$B_3714_out0[3:3];
assign v$_3482_out0 = { v$G15_2300_out0,v$G16_1803_out0 };
assign v$_3483_out0 = { v$G15_2301_out0,v$G16_1804_out0 };
assign v$C5_3633_out0 = v$SEL22_960_out0;
assign v$C1_3693_out0 = v$SEL21_756_out0;
assign v$SEL13_3870_out0 = v$B_3712_out0[2:2];
assign v$SEL13_3871_out0 = v$B_3713_out0[2:2];
assign v$SEL13_3872_out0 = v$B_3714_out0[2:2];
assign v$SEL16_3938_out0 = v$B_3712_out0[8:8];
assign v$SEL16_3939_out0 = v$B_3713_out0[8:8];
assign v$SEL16_3940_out0 = v$B_3714_out0[8:8];
assign v$SEL23_3969_out0 = v$C_3602_out0[6:6];
assign v$SEL23_3971_out0 = v$C_3604_out0[6:6];
assign v$C2_3991_out0 = v$SEL25_4657_out0;
assign v$SEL5_4030_out0 = v$A_3705_out0[8:8];
assign v$SEL5_4031_out0 = v$A_3706_out0[8:8];
assign v$SEL5_4032_out0 = v$A_3707_out0[8:8];
assign v$SEL5_4148_out0 = v$A_3570_out0[5:5];
assign v$SEL21_4310_out0 = v$C_4519_out0[6:6];
assign v$SEL17_4472_out0 = v$B_3712_out0[7:7];
assign v$SEL17_4473_out0 = v$B_3713_out0[7:7];
assign v$SEL17_4474_out0 = v$B_3714_out0[7:7];
assign v$SEL20_4544_out0 = v$C_3602_out0[0:0];
assign v$SEL20_4546_out0 = v$C_3604_out0[0:0];
assign v$SEL28_4556_out0 = v$A_3570_out0[9:9];
assign v$SEL25_4656_out0 = v$C_3602_out0[2:2];
assign v$SEL25_4658_out0 = v$C_3604_out0[2:2];
assign v$SEL25_4721_out0 = v$C_4519_out0[2:2];
assign v$SEL8_4726_out0 = v$A_3705_out0[7:7];
assign v$SEL8_4727_out0 = v$A_3706_out0[7:7];
assign v$SEL8_4728_out0 = v$A_3707_out0[7:7];
assign v$C3_4734_out0 = v$SEL24_1793_out0;
assign v$SEL10_4866_out0 = v$C_4519_out0[8:8];
assign v$C8_4925_out0 = v$SEL26_1708_out0;
assign v$SEL7_5192_out0 = v$A_3705_out0[3:3];
assign v$SEL7_5193_out0 = v$A_3706_out0[3:3];
assign v$SEL7_5194_out0 = v$A_3707_out0[3:3];
assign v$Toshift_5200_out0 = v$SHIFTSIGNIFICANT_5041_out0;
assign v$SEL14_5216_out0 = v$C_4519_out0[7:7];
assign v$G5_5360_out0 = v$A_4971_out0 && v$B_61_out0;
assign v$G5_5365_out0 = v$A_4976_out0 && v$B_66_out0;
assign v$G5_5366_out0 = v$A_4977_out0 && v$B_67_out0;
assign v$G5_5371_out0 = v$A_4982_out0 && v$B_72_out0;
assign v$G5_5372_out0 = v$A_4983_out0 && v$B_73_out0;
assign v$G5_5376_out0 = v$A_4987_out0 && v$B_77_out0;
assign v$C0_5421_out0 = v$SEL20_4545_out0;
assign v$C3_29_out0 = v$SEL11_3136_out0;
assign v$A5_51_out0 = v$SEL6_1042_out0;
assign v$A5_52_out0 = v$SEL6_1043_out0;
assign v$A5_53_out0 = v$SEL6_1044_out0;
assign v$C2_199_out0 = v$SEL25_4721_out0;
assign v$A6_211_out0 = v$SEL2_605_out0;
assign v$A2_313_out0 = v$SEL4_3162_out0;
assign v$A2_314_out0 = v$SEL4_3163_out0;
assign v$A2_315_out0 = v$SEL4_3164_out0;
assign v$A3_370_out0 = v$SEL27_919_out0;
assign v$A0_551_out0 = v$SEL9_3387_out0;
assign v$A0_552_out0 = v$SEL9_3388_out0;
assign v$A0_553_out0 = v$SEL9_3389_out0;
assign v$C_639_out0 = v$G5_5360_out0;
assign v$C_644_out0 = v$G5_5365_out0;
assign v$C_645_out0 = v$G5_5366_out0;
assign v$C_650_out0 = v$G5_5371_out0;
assign v$C_651_out0 = v$G5_5372_out0;
assign v$C_655_out0 = v$G5_5376_out0;
assign v$C9_699_out0 = v$SEL30_1615_out0;
assign v$A1_732_out0 = v$SEL1_3306_out0;
assign v$A1_733_out0 = v$SEL1_3307_out0;
assign v$A1_734_out0 = v$SEL1_3308_out0;
assign v$B2_765_out0 = v$SEL13_3870_out0;
assign v$B2_766_out0 = v$SEL13_3871_out0;
assign v$B2_767_out0 = v$SEL13_3872_out0;
assign v$A0_915_out0 = v$SEL17_994_out0;
assign v$A3_1053_out0 = v$SEL7_5192_out0;
assign v$A3_1054_out0 = v$SEL7_5193_out0;
assign v$A3_1055_out0 = v$SEL7_5194_out0;
assign v$C0_1109_out0 = v$SEL24_1409_out0;
assign v$A9_1282_out0 = v$SEL28_4556_out0;
assign v$C1_1392_out0 = v$SEL3_1664_out0;
assign v$A8_1454_out0 = v$SEL22_2924_out0;
assign v$A8_1557_out0 = v$SEL5_4030_out0;
assign v$A8_1558_out0 = v$SEL5_4031_out0;
assign v$A8_1559_out0 = v$SEL5_4032_out0;
assign v$B4_1868_out0 = v$SEL10_1159_out0;
assign v$B4_1869_out0 = v$SEL10_1160_out0;
assign v$B4_1870_out0 = v$SEL10_1161_out0;
assign v$G0_1975_out0 = v$A_4971_out0 && v$G4_1331_out0;
assign v$G0_1980_out0 = v$A_4976_out0 && v$G4_1336_out0;
assign v$G0_1981_out0 = v$A_4977_out0 && v$G4_1337_out0;
assign v$G0_1986_out0 = v$A_4982_out0 && v$G4_1342_out0;
assign v$G0_1987_out0 = v$A_4983_out0 && v$G4_1343_out0;
assign v$G0_1991_out0 = v$A_4987_out0 && v$G4_1347_out0;
assign v$B7_2161_out0 = v$SEL17_4472_out0;
assign v$B7_2162_out0 = v$SEL17_4473_out0;
assign v$B7_2163_out0 = v$SEL17_4474_out0;
assign v$B8_2202_out0 = v$SEL16_3938_out0;
assign v$B8_2203_out0 = v$SEL16_3939_out0;
assign v$B8_2204_out0 = v$SEL16_3940_out0;
assign v$A4_2222_out0 = v$SEL1_3203_out0;
assign v$C7_2318_out0 = v$SEL27_2608_out0;
assign v$C7_2320_out0 = v$SEL27_2610_out0;
assign v$A4_2443_out0 = v$SEL3_358_out0;
assign v$A4_2444_out0 = v$SEL3_359_out0;
assign v$A4_2445_out0 = v$SEL3_360_out0;
assign v$C8_2450_out0 = v$SEL10_4866_out0;
assign v$G1_2518_out0 = v$G3_2803_out0 && v$B_61_out0;
assign v$G1_2524_out0 = v$G3_2809_out0 && v$B_67_out0;
assign v$G1_2529_out0 = v$G3_2814_out0 && v$B_72_out0;
assign v$G1_2530_out0 = v$G3_2815_out0 && v$B_73_out0;
assign v$G1_2534_out0 = v$G3_2819_out0 && v$B_77_out0;
assign v$XOR1_2651_out0 = v$Toshift_5200_out0 ^ v$MUX1_4000_out0;
assign v$C6_2675_out0 = v$SEL23_3969_out0;
assign v$C6_2677_out0 = v$SEL23_3971_out0;
assign v$A2_2730_out0 = v$SEL15_832_out0;
assign v$B5_3028_out0 = v$SEL12_2082_out0;
assign v$B5_3029_out0 = v$SEL12_2083_out0;
assign v$B5_3030_out0 = v$SEL12_2084_out0;
assign v$C4_3419_out0 = v$SEL19_1487_out0;
assign v$C4_3421_out0 = v$SEL19_1489_out0;
assign v$C5_3632_out0 = v$SEL22_959_out0;
assign v$C5_3634_out0 = v$SEL22_961_out0;
assign v$C1_3692_out0 = v$SEL21_755_out0;
assign v$C1_3694_out0 = v$SEL21_757_out0;
assign v$A6_3769_out0 = v$SEL2_740_out0;
assign v$A6_3770_out0 = v$SEL2_741_out0;
assign v$A6_3771_out0 = v$SEL2_742_out0;
assign v$A1_3822_out0 = v$SEL16_1897_out0;
assign v$C2_3990_out0 = v$SEL25_4656_out0;
assign v$C2_3992_out0 = v$SEL25_4658_out0;
assign v$A7_4165_out0 = v$SEL26_1765_out0;
assign v$C4_4230_out0 = v$SEL8_1505_out0;
assign v$C7_4234_out0 = v$SEL14_5216_out0;
assign v$A7_4560_out0 = v$SEL8_4726_out0;
assign v$A7_4561_out0 = v$SEL8_4727_out0;
assign v$A7_4562_out0 = v$SEL8_4728_out0;
assign v$C5_4631_out0 = v$SEL4_40_out0;
assign v$C3_4733_out0 = v$SEL24_1792_out0;
assign v$C3_4735_out0 = v$SEL24_1794_out0;
assign v$A5_4740_out0 = v$SEL5_4148_out0;
assign v$B6_4851_out0 = v$SEL11_2550_out0;
assign v$B6_4852_out0 = v$SEL11_2551_out0;
assign v$B6_4853_out0 = v$SEL11_2552_out0;
assign v$C8_4924_out0 = v$SEL26_1707_out0;
assign v$C8_4926_out0 = v$SEL26_1709_out0;
assign v$B3_5123_out0 = v$SEL18_3450_out0;
assign v$B3_5124_out0 = v$SEL18_3451_out0;
assign v$B3_5125_out0 = v$SEL18_3452_out0;
assign v$C6_5172_out0 = v$SEL21_4310_out0;
assign v$_5276_out0 = { v$_3547_out0,v$_3482_out0 };
assign v$_5277_out0 = { v$_3548_out0,v$_3483_out0 };
assign v$B0_5314_out0 = v$SEL15_1364_out0;
assign v$B0_5315_out0 = v$SEL15_1365_out0;
assign v$B0_5316_out0 = v$SEL15_1366_out0;
assign v$B1_5323_out0 = v$SEL14_1492_out0;
assign v$B1_5324_out0 = v$SEL14_1493_out0;
assign v$B1_5325_out0 = v$SEL14_1494_out0;
assign v$C0_5420_out0 = v$SEL20_4544_out0;
assign v$C0_5422_out0 = v$SEL20_4546_out0;
assign v$G2_430_out0 = v$G0_1975_out0 || v$G1_2518_out0;
assign v$G2_435_out0 = v$G0_1980_out0 || v$G1_2523_out0;
assign v$G2_436_out0 = v$G0_1981_out0 || v$G1_2524_out0;
assign v$G2_441_out0 = v$G0_1986_out0 || v$G1_2529_out0;
assign v$G2_442_out0 = v$G0_1987_out0 || v$G1_2530_out0;
assign v$G2_446_out0 = v$G0_1991_out0 || v$G1_2534_out0;
assign {v$A4_520_out1,v$A4_520_out0 } = v$B4_1868_out0 + v$C4_3419_out0 + v$A4_2443_out0;
assign {v$A4_521_out1,v$A4_521_out0 } = v$B4_1869_out0 + v$C4_3420_out0 + v$A4_2444_out0;
assign {v$A4_522_out1,v$A4_522_out0 } = v$B4_1870_out0 + v$C4_3421_out0 + v$A4_2445_out0;
assign v$_836_out0 = { v$C2_3555_out0,v$C_639_out0 };
assign {v$A6_1091_out1,v$A6_1091_out0 } = v$B3_5123_out0 + v$C3_4733_out0 + v$A3_1053_out0;
assign {v$A6_1092_out1,v$A6_1092_out0 } = v$B3_5124_out0 + v$C3_4734_out0 + v$A3_1054_out0;
assign {v$A6_1093_out1,v$A6_1093_out0 } = v$B3_5125_out0 + v$C3_4735_out0 + v$A3_1055_out0;
assign v$_1386_out0 = { v$C1_4681_out0,v$C_644_out0 };
assign {v$A7_1863_out1,v$A7_1863_out0 } = v$B7_2161_out0 + v$C7_2318_out0 + v$A7_4560_out0;
assign {v$A7_1864_out1,v$A7_1864_out0 } = v$B7_2162_out0 + v$C7_2319_out0 + v$A7_4561_out0;
assign {v$A7_1865_out1,v$A7_1865_out0 } = v$B7_2163_out0 + v$C7_2320_out0 + v$A7_4562_out0;
assign {v$A2_2603_out1,v$A2_2603_out0 } = v$B1_5323_out0 + v$C1_3692_out0 + v$A1_732_out0;
assign {v$A2_2604_out1,v$A2_2604_out0 } = v$B1_5324_out0 + v$C1_3693_out0 + v$A1_733_out0;
assign {v$A2_2605_out1,v$A2_2605_out0 } = v$B1_5325_out0 + v$C1_3694_out0 + v$A1_734_out0;
assign {v$A3_2872_out1,v$A3_2872_out0 } = v$B2_765_out0 + v$C2_3990_out0 + v$A2_313_out0;
assign {v$A3_2873_out1,v$A3_2873_out0 } = v$B2_766_out0 + v$C2_3991_out0 + v$A2_314_out0;
assign {v$A3_2874_out1,v$A3_2874_out0 } = v$B2_767_out0 + v$C2_3992_out0 + v$A2_315_out0;
assign v$_3078_out0 = { v$C4_1537_out0,v$C_655_out0 };
assign {v$A1_3679_out1,v$A1_3679_out0 } = v$_4828_out0 + v$XOR1_2651_out0 + v$SUB_4899_out0;
assign {v$A8_3701_out1,v$A8_3701_out0 } = v$B6_4851_out0 + v$C6_2675_out0 + v$A6_3769_out0;
assign {v$A8_3702_out1,v$A8_3702_out0 } = v$B6_4852_out0 + v$C6_2676_out0 + v$A6_3770_out0;
assign {v$A8_3703_out1,v$A8_3703_out0 } = v$B6_4853_out0 + v$C6_2677_out0 + v$A6_3771_out0;
assign {v$A1_3716_out1,v$A1_3716_out0 } = v$B0_5314_out0 + v$C0_5420_out0 + v$A0_551_out0;
assign {v$A1_3717_out1,v$A1_3717_out0 } = v$B0_5315_out0 + v$C0_5421_out0 + v$A0_552_out0;
assign {v$A1_3718_out1,v$A1_3718_out0 } = v$B0_5316_out0 + v$C0_5422_out0 + v$A0_553_out0;
assign v$_3924_out0 = { v$_3591_out0,v$_5276_out0 };
assign v$_3925_out0 = { v$_3592_out0,v$_5277_out0 };
assign {v$A9_4400_out1,v$A9_4400_out0 } = v$B8_2202_out0 + v$C8_4924_out0 + v$A8_1557_out0;
assign {v$A9_4401_out1,v$A9_4401_out0 } = v$B8_2203_out0 + v$C8_4925_out0 + v$A8_1558_out0;
assign {v$A9_4402_out1,v$A9_4402_out0 } = v$B8_2204_out0 + v$C8_4926_out0 + v$A8_1559_out0;
assign {v$A5_5012_out1,v$A5_5012_out0 } = v$B5_3028_out0 + v$C5_3632_out0 + v$A5_51_out0;
assign {v$A5_5013_out1,v$A5_5013_out0 } = v$B5_3029_out0 + v$C5_3633_out0 + v$A5_52_out0;
assign {v$A5_5014_out1,v$A5_5014_out0 } = v$B5_3030_out0 + v$C5_3634_out0 + v$A5_53_out0;
assign v$S01_192_out0 = v$A2_2603_out0;
assign v$S01_193_out0 = v$A2_2604_out0;
assign v$S01_194_out0 = v$A2_2605_out0;
assign v$S15_459_out0 = v$A5_5012_out1;
assign v$S15_460_out0 = v$A5_5013_out1;
assign v$S15_461_out0 = v$A5_5014_out1;
assign v$S04_928_out0 = v$A4_520_out0;
assign v$S04_929_out0 = v$A4_521_out0;
assign v$S04_930_out0 = v$A4_522_out0;
assign v$S02_1073_out0 = v$A3_2872_out0;
assign v$S02_1074_out0 = v$A3_2873_out0;
assign v$S02_1075_out0 = v$A3_2874_out0;
assign v$S00_1129_out0 = v$A1_3716_out0;
assign v$S00_1130_out0 = v$A1_3717_out0;
assign v$S00_1131_out0 = v$A1_3718_out0;
assign v$S07_1255_out0 = v$A7_1863_out0;
assign v$S07_1256_out0 = v$A7_1864_out0;
assign v$S07_1257_out0 = v$A7_1865_out0;
assign v$S18_1962_out0 = v$A9_4400_out1;
assign v$S18_1963_out0 = v$A9_4401_out1;
assign v$S18_1964_out0 = v$A9_4402_out1;
assign v$S11_2562_out0 = v$A2_2603_out1;
assign v$S11_2563_out0 = v$A2_2604_out1;
assign v$S11_2564_out0 = v$A2_2605_out1;
assign v$S17_2862_out0 = v$A7_1863_out1;
assign v$S17_2863_out0 = v$A7_1864_out1;
assign v$S17_2864_out0 = v$A7_1865_out1;
assign v$S05_2989_out0 = v$A5_5012_out0;
assign v$S05_2990_out0 = v$A5_5013_out0;
assign v$S05_2991_out0 = v$A5_5014_out0;
assign v$S03_3015_out0 = v$A6_1091_out0;
assign v$S03_3016_out0 = v$A6_1092_out0;
assign v$S03_3017_out0 = v$A6_1093_out0;
assign v$_3101_out0 = { v$_745_out0,v$_3924_out0 };
assign v$_3102_out0 = { v$_746_out0,v$_3925_out0 };
assign v$S14_3380_out0 = v$A4_520_out1;
assign v$S14_3381_out0 = v$A4_521_out1;
assign v$S14_3382_out0 = v$A4_522_out1;
assign v$S13_3437_out0 = v$A6_1091_out1;
assign v$S13_3438_out0 = v$A6_1092_out1;
assign v$S13_3439_out0 = v$A6_1093_out1;
assign v$S10_3472_out0 = v$A1_3716_out1;
assign v$S10_3473_out0 = v$A1_3717_out1;
assign v$S10_3474_out0 = v$A1_3718_out1;
assign v$COUT_4071_out0 = v$A1_3679_out1;
assign v$S_4176_out0 = v$G2_430_out0;
assign v$S_4181_out0 = v$G2_435_out0;
assign v$S_4182_out0 = v$G2_436_out0;
assign v$S_4187_out0 = v$G2_441_out0;
assign v$S_4188_out0 = v$G2_442_out0;
assign v$S_4192_out0 = v$G2_446_out0;
assign v$S06_4368_out0 = v$A8_3701_out0;
assign v$S06_4369_out0 = v$A8_3702_out0;
assign v$S06_4370_out0 = v$A8_3703_out0;
assign v$S12_4799_out0 = v$A3_2872_out1;
assign v$S12_4800_out0 = v$A3_2873_out1;
assign v$S12_4801_out0 = v$A3_2874_out1;
assign v$S16_4892_out0 = v$A8_3701_out1;
assign v$S16_4893_out0 = v$A8_3702_out1;
assign v$S16_4894_out0 = v$A8_3703_out1;
assign v$SUM_5158_out0 = v$A1_3679_out0;
assign v$S08_5272_out0 = v$A9_4400_out0;
assign v$S08_5273_out0 = v$A9_4401_out0;
assign v$S08_5274_out0 = v$A9_4402_out0;
assign v$_840_out0 = { v$S10_3472_out0,v$S11_2562_out0 };
assign v$_841_out0 = { v$S10_3473_out0,v$S11_2563_out0 };
assign v$_842_out0 = { v$S10_3474_out0,v$S11_2564_out0 };
assign v$_1431_out0 = { v$S04_928_out0,v$S05_2989_out0 };
assign v$_1432_out0 = { v$S04_929_out0,v$S05_2990_out0 };
assign v$_1433_out0 = { v$S04_930_out0,v$S05_2991_out0 };
assign v$_1562_out0 = { v$SEL1_4808_out0,v$S_4181_out0 };
assign v$_1608_out0 = { v$S02_1073_out0,v$S03_3015_out0 };
assign v$_1609_out0 = { v$S02_1074_out0,v$S03_3016_out0 };
assign v$_1610_out0 = { v$S02_1075_out0,v$S03_3017_out0 };
assign v$_1809_out0 = { v$S_4187_out0,v$SEL21_2848_out0 };
assign v$_2354_out0 = { v$S12_4799_out0,v$S13_3437_out0 };
assign v$_2355_out0 = { v$S12_4800_out0,v$S13_3438_out0 };
assign v$_2356_out0 = { v$S12_4801_out0,v$S13_3439_out0 };
assign v$_2978_out0 = { v$S16_4892_out0,v$S17_2862_out0 };
assign v$_2979_out0 = { v$S16_4893_out0,v$S17_2863_out0 };
assign v$_2980_out0 = { v$S16_4894_out0,v$S17_2864_out0 };
assign v$_3066_out0 = { v$_272_out0,v$S_4176_out0 };
assign v$_3364_out0 = { v$S_4188_out0,v$SEL33_1822_out0 };
assign v$_3625_out0 = { v$S06_4368_out0,v$S07_1255_out0 };
assign v$_3626_out0 = { v$S06_4369_out0,v$S07_1256_out0 };
assign v$_3627_out0 = { v$S06_4370_out0,v$S07_1257_out0 };
assign v$_3638_out0 = { v$S00_1129_out0,v$S01_192_out0 };
assign v$_3639_out0 = { v$S00_1130_out0,v$S01_193_out0 };
assign v$_3640_out0 = { v$S00_1131_out0,v$S01_194_out0 };
assign v$_3667_out0 = v$SUM_5158_out0[0:0];
assign v$_3667_out1 = v$SUM_5158_out0[12:12];
assign v$_3847_out0 = { v$_5429_out0,v$S_4192_out0 };
assign v$G1_4094_out0 = v$COUT_4071_out0 && v$G2_4803_out0;
assign v$_4127_out0 = { v$S14_3380_out0,v$S15_459_out0 };
assign v$_4128_out0 = { v$S14_3381_out0,v$S15_460_out0 };
assign v$_4129_out0 = { v$S14_3382_out0,v$S15_461_out0 };
assign v$X_4521_out0 = v$_3101_out0;
assign v$X_4522_out0 = v$_3102_out0;
assign v$_4858_out0 = { v$S_4182_out0,v$SEL26_529_out0 };
assign v$_1604_out0 = { v$_4127_out0,v$_2978_out0 };
assign v$_1605_out0 = { v$_4128_out0,v$_2979_out0 };
assign v$_1606_out0 = { v$_4129_out0,v$_2980_out0 };
assign v$STICKY_1727_out0 = v$_3667_out0;
assign v$_2659_out0 = { v$_1431_out0,v$_3625_out0 };
assign v$_2660_out0 = { v$_1432_out0,v$_3626_out0 };
assign v$_2661_out0 = { v$_1433_out0,v$_3627_out0 };
assign v$ANDOUT_3462_out0 = v$X_4521_out0;
assign v$ANDOUT_3463_out0 = v$X_4522_out0;
assign v$_4158_out0 = { v$_3638_out0,v$_1608_out0 };
assign v$_4159_out0 = { v$_3639_out0,v$_1609_out0 };
assign v$_4160_out0 = { v$_3640_out0,v$_1610_out0 };
assign v$_4754_out0 = { v$_840_out0,v$_2354_out0 };
assign v$_4755_out0 = { v$_841_out0,v$_2355_out0 };
assign v$_4756_out0 = { v$_842_out0,v$_2356_out0 };
assign v$DETECT1_5247_out0 = v$G1_4094_out0;
assign v$MUX6_796_out0 = v$G12_5243_out0 ? v$ANDOUT_3462_out0 : v$MUX4_5267_out0;
assign v$MUX6_797_out0 = v$G12_5244_out0 ? v$ANDOUT_3463_out0 : v$MUX4_5268_out0;
assign v$_2463_out0 = { v$_2659_out0,v$S08_5272_out0 };
assign v$_2464_out0 = { v$_2660_out0,v$S08_5273_out0 };
assign v$_2465_out0 = { v$_2661_out0,v$S08_5274_out0 };
assign v$G3_2968_out0 = v$EQ1_4746_out0 && v$DETECT1_5247_out0;
assign v$_4323_out0 = { v$_1604_out0,v$S18_1962_out0 };
assign v$_4324_out0 = { v$_1605_out0,v$S18_1963_out0 };
assign v$_4325_out0 = { v$_1606_out0,v$S18_1964_out0 };
assign v$DETECT1_4467_out0 = v$DETECT1_5247_out0;
assign v$_5254_out0 = { v$_3667_out1,v$DETECT1_5247_out0 };
assign v$_217_out0 = { v$_4754_out0,v$_4323_out0 };
assign v$_218_out0 = { v$_4755_out0,v$_4324_out0 };
assign v$_219_out0 = { v$_4756_out0,v$_4325_out0 };
assign v$ALUOUT_1768_out0 = v$MUX6_796_out0;
assign v$ALUOUT_1769_out0 = v$MUX6_797_out0;
assign v$DETECT1_2843_out0 = v$DETECT1_4467_out0;
assign v$OVERFLOW_2960_out0 = v$G3_2968_out0;
assign v$_3865_out0 = { v$_4158_out0,v$_2463_out0 };
assign v$_3866_out0 = { v$_4159_out0,v$_2464_out0 };
assign v$_3867_out0 = { v$_4160_out0,v$_2465_out0 };
assign v$ADD2_4212_out0 = v$_5254_out0;
assign v$ALUOUT_545_out0 = v$ALUOUT_1768_out0;
assign v$ALUOUT_546_out0 = v$ALUOUT_1769_out0;
assign v$S0_1260_out0 = v$_3865_out0;
assign v$S0_1261_out0 = v$_3866_out0;
assign v$S0_1262_out0 = v$_3867_out0;
assign v$MUX2_1808_out0 = v$DETECT1_5247_out0 ? v$ADD2_4212_out0 : v$SUM_5158_out0;
assign v$DETECT1_1926_out0 = v$DETECT1_2843_out0;
assign v$S1_4225_out0 = v$_217_out0;
assign v$S1_4226_out0 = v$_218_out0;
assign v$S1_4227_out0 = v$_219_out0;
assign v$G2_5351_out0 = v$G1_706_out0 || v$OVERFLOW_2960_out0;
assign v$_196_out0 = { v$_1562_out0,v$S0_1261_out0 };
assign v$_222_out0 = { v$_3066_out0,v$S0_1260_out0 };
assign v$EXCEPTION_855_out0 = v$G2_5351_out0;
assign v$_1825_out0 = { v$S1_4227_out0,v$C_651_out0 };
assign v$_2500_out0 = { v$S1_4225_out0,v$C_645_out0 };
assign v$MUX1_3564_out0 = v$IR15_322_out0 ? v$ALUOUT_545_out0 : v$REGDIN_1934_out0;
assign v$MUX1_3565_out0 = v$IR15_323_out0 ? v$ALUOUT_546_out0 : v$REGDIN_1935_out0;
assign v$ALUOUT_3587_out0 = v$ALUOUT_545_out0;
assign v$ALUOUT_3588_out0 = v$ALUOUT_546_out0;
assign v$ALUOUT_3789_out0 = v$ALUOUT_545_out0;
assign v$ALUOUT_3790_out0 = v$ALUOUT_546_out0;
assign v$_4319_out0 = { v$S1_4226_out0,v$C_650_out0 };
assign v$OUTPUT_4621_out0 = v$MUX2_1808_out0;
assign v$_4747_out0 = { v$_3847_out0,v$S0_1262_out0 };
assign v$_771_out0 = { v$_1386_out0,v$_4319_out0 };
assign v$_1371_out0 = { v$_3078_out0,v$_1825_out0 };
assign v$IN_1445_out0 = v$OUTPUT_4621_out0;
assign v$ALUOUT_1496_out0 = v$ALUOUT_3587_out0;
assign v$ALUOUT_1497_out0 = v$ALUOUT_3588_out0;
assign v$_1536_out0 = { v$_836_out0,v$_2500_out0 };
assign v$INPUT_3073_out0 = v$OUTPUT_4621_out0;
assign v$DIN3_3861_out0 = v$MUX1_3564_out0;
assign v$DIN3_3862_out0 = v$MUX1_3565_out0;
assign v$_4532_out0 = { v$_4747_out0,v$_3364_out0 };
assign v$_4564_out0 = { v$_222_out0,v$_4858_out0 };
assign v$_4638_out0 = { v$_196_out0,v$_1809_out0 };
assign v$ALUOUT_5256_out0 = v$ALUOUT_3789_out0;
assign v$ALUOUT_5257_out0 = v$ALUOUT_3790_out0;
assign v$EXCEPTION_5275_out0 = v$EXCEPTION_855_out0;
assign v$SEL18_26_out0 = v$INPUT_3073_out0[3:3];
assign v$MUX12_152_out0 = v$RET_2085_out0 ? v$R1S_279_out0 : v$DIN3_3861_out0;
assign v$MUX12_153_out0 = v$RET_2086_out0 ? v$R1S_280_out0 : v$DIN3_3862_out0;
assign v$SEL5_267_out0 = v$INPUT_3073_out0[10:10];
assign v$SEL15_469_out0 = v$INPUT_3073_out0[4:4];
assign v$SEL14_1155_out0 = v$INPUT_3073_out0[7:7];
assign v$SEL12_1174_out0 = v$INPUT_3073_out0[12:12];
assign v$MUX11_1403_out0 = v$RET_2085_out0 ? v$R0S_1142_out0 : v$DIN3_3861_out0;
assign v$MUX11_1404_out0 = v$RET_2086_out0 ? v$R0S_1143_out0 : v$DIN3_3862_out0;
assign v$SEL7_1406_out0 = v$INPUT_3073_out0[8:8];
assign v$SEL6_1561_out0 = v$INPUT_3073_out0[9:9];
assign v$L5_1655_out0 = v$_1371_out0;
assign v$MUX14_1674_out0 = v$RET_2085_out0 ? v$R3S_4764_out0 : v$DIN3_3861_out0;
assign v$MUX14_1675_out0 = v$RET_2086_out0 ? v$R3S_4765_out0 : v$DIN3_3862_out0;
assign v$SEL21_2093_out0 = v$INPUT_3073_out0[0:0];
assign v$L1_2240_out0 = v$_771_out0;
assign v$SEL20_2272_out0 = v$INPUT_3073_out0[1:1];
assign v$L0_2414_out0 = v$_4638_out0;
assign v$L2_3025_out0 = v$_4564_out0;
assign v$INPUT_3065_out0 = v$IN_1445_out0;
assign v$SEL13_3457_out0 = v$INPUT_3073_out0[6:6];
assign v$SEL17_3946_out0 = v$INPUT_3073_out0[2:2];
assign v$SEL16_4040_out0 = v$INPUT_3073_out0[5:5];
assign v$MUX13_4054_out0 = v$RET_2085_out0 ? v$R2S_1379_out0 : v$DIN3_3861_out0;
assign v$MUX13_4055_out0 = v$RET_2086_out0 ? v$R2S_1380_out0 : v$DIN3_3862_out0;
assign v$SEL1_4768_out0 = v$INPUT_3073_out0[11:11];
assign v$L3_5181_out0 = v$_1536_out0;
assign v$L4_5246_out0 = v$_4532_out0;
assign v$SEL45_173_out0 = v$L0_2414_out0[12:3];
assign v$G52_303_out0 = ! v$SEL15_469_out0;
assign v$G66_558_out0 = ! v$SEL21_2093_out0;
assign v$G46_561_out0 = ! v$SEL13_3457_out0;
assign v$SEL50_736_out0 = v$L4_5246_out0[6:6];
assign v$SEL55_752_out0 = v$L3_5181_out0[5:5];
assign v$G19_787_out0 = ! v$SEL5_267_out0;
assign v$SEL52_902_out0 = v$L5_1655_out0[15:8];
assign v$SEL46_1049_out0 = v$L1_2240_out0[2:2];
assign v$G17_1083_out0 = ! v$SEL1_4768_out0;
assign v$SEL43_1228_out0 = v$L1_2240_out0[12:3];
assign v$G39_1319_out0 = ! v$SEL12_1174_out0;
assign v$SEL56_1474_out0 = v$L4_5246_out0[7:7];
assign v$SEL66_1553_out0 = v$L5_1655_out0[17:17];
assign v$SEL64_2195_out0 = v$L5_1655_out0[18:18];
assign v$G40_2290_out0 = ! v$SEL7_1406_out0;
assign v$SEL51_2334_out0 = v$L4_5246_out0[15:8];
assign v$G45_2793_out0 = ! v$SEL14_1155_out0;
assign v$SEL41_2794_out0 = v$L2_3025_out0[12:3];
assign v$SEL90_2866_out0 = v$L2_3025_out0[13:13];
assign v$SEL57_2938_out0 = v$L3_5181_out0[7:7];
assign v$SEL49_3044_out0 = v$L3_5181_out0[15:8];
assign v$G22_3337_out0 = ! v$SEL6_1561_out0;
assign v$G51_3597_out0 = ! v$SEL16_4040_out0;
assign v$SEL65_3615_out0 = v$L5_1655_out0[16:16];
assign v$SEL42_3888_out0 = v$L0_2414_out0[2:2];
assign v$SEL63_3931_out0 = v$L4_5246_out0[18:18];
assign v$SEL53_4486_out0 = v$L3_5181_out0[6:6];
assign v$SEL47_4498_out0 = v$L2_3025_out0[15:14];
assign v$SEL58_4499_out0 = v$L4_5246_out0[16:16];
assign v$G58_4585_out0 = ! v$SEL17_3946_out0;
assign v$SEL59_4818_out0 = v$L4_5246_out0[17:17];
assign v$SEL48_4857_out0 = v$L0_2414_out0[1:0];
assign v$G57_4885_out0 = ! v$SEL18_26_out0;
assign v$G62_4943_out0 = ! v$SEL20_2272_out0;
assign v$12_5203_out0 = v$SEL12_1174_out0;
assign v$B_62_out0 = v$SEL63_3931_out0;
assign v$B_68_out0 = v$SEL50_736_out0;
assign v$B_69_out0 = v$SEL46_1049_out0;
assign v$B_71_out0 = v$SEL56_1474_out0;
assign v$B_74_out0 = v$SEL58_4499_out0;
assign v$B_75_out0 = v$SEL59_4818_out0;
assign v$MUX13_850_out0 = v$12_5203_out0 ? v$C2_4460_out0 : v$C1_2299_out0;
assign v$G18_2014_out0 = v$G17_1083_out0 && v$G39_1319_out0;
assign v$B_2057_out0 = v$SEL51_2334_out0;
assign v$C_2732_out0 = v$SEL49_3044_out0;
assign v$G6_3368_out0 = v$SEL1_4768_out0 && v$G39_1319_out0;
assign v$A_3569_out0 = v$SEL43_1228_out0;
assign v$B_3841_out0 = v$SEL45_173_out0;
assign v$C_4518_out0 = v$SEL41_2794_out0;
assign v$A_4699_out0 = v$SEL52_902_out0;
assign v$A_4972_out0 = v$SEL64_2195_out0;
assign v$A_4978_out0 = v$SEL53_4486_out0;
assign v$A_4979_out0 = v$SEL42_3888_out0;
assign v$A_4981_out0 = v$SEL57_2938_out0;
assign v$A_4984_out0 = v$SEL65_3615_out0;
assign v$A_4985_out0 = v$SEL66_1553_out0;
assign v$_5278_out0 = { v$C8_13_out0,v$SEL55_752_out0 };
assign v$SEL23_9_out0 = v$B_2057_out0[7:7];
assign v$SEL4_39_out0 = v$C_4518_out0[5:5];
assign v$SEL29_97_out0 = v$B_3841_out0[9:9];
assign v$G20_319_out0 = v$SEL5_267_out0 && v$G18_2014_out0;
assign v$SEL8_355_out0 = v$C_2732_out0[4:4];
assign v$SEL27_412_out0 = v$A_4699_out0[3:3];
assign v$SEL15_496_out0 = v$A_4699_out0[2:2];
assign v$SEL23_585_out0 = v$B_3841_out0[7:7];
assign v$SEL2_604_out0 = v$A_3569_out0[6:6];
assign v$SEL4_768_out0 = v$C_2732_out0[5:5];
assign v$SEL15_831_out0 = v$A_3569_out0[2:2];
assign v$SEL27_918_out0 = v$A_3569_out0[3:3];
assign v$SEL21_969_out0 = v$C_2732_out0[6:6];
assign v$SEL17_993_out0 = v$A_3569_out0[0:0];
assign v$SEL19_1071_out0 = v$B_2057_out0[2:2];
assign v$SEL3_1276_out0 = v$C_2732_out0[1:1];
assign v$SEL1_1279_out0 = v$A_4699_out0[4:4];
assign v$G4_1332_out0 = ! v$B_62_out0;
assign v$G4_1338_out0 = ! v$B_68_out0;
assign v$G4_1339_out0 = ! v$B_69_out0;
assign v$G4_1341_out0 = ! v$B_71_out0;
assign v$G4_1344_out0 = ! v$B_74_out0;
assign v$G4_1345_out0 = ! v$B_75_out0;
assign v$SEL24_1408_out0 = v$C_4518_out0[0:0];
assign v$G23_1485_out0 = v$G19_787_out0 && v$G18_2014_out0;
assign v$SEL8_1504_out0 = v$C_4518_out0[4:4];
assign v$SEL6_1508_out0 = v$B_3841_out0[4:4];
assign v$SEL19_1533_out0 = v$B_3841_out0[2:2];
assign v$SEL30_1614_out0 = v$C_4518_out0[9:9];
assign v$SEL3_1663_out0 = v$C_4518_out0[1:1];
assign v$SEL25_1731_out0 = v$C_2732_out0[2:2];
assign v$SEL26_1764_out0 = v$A_3569_out0[7:7];
assign v$SEL20_1842_out0 = v$B_3841_out0[8:8];
assign v$SEL7_1848_out0 = v$B_3841_out0[0:0];
assign v$SEL16_1896_out0 = v$A_3569_out0[1:1];
assign v$SEL16_2266_out0 = v$A_4699_out0[1:1];
assign v$SEL18_2406_out0 = v$B_2057_out0[3:3];
assign v$SEL12_2598_out0 = v$B_2057_out0[5:5];
assign v$SEL6_2599_out0 = v$B_2057_out0[4:4];
assign v$G3_2804_out0 = ! v$A_4972_out0;
assign v$G3_2810_out0 = ! v$A_4978_out0;
assign v$G3_2811_out0 = ! v$A_4979_out0;
assign v$G3_2813_out0 = ! v$A_4981_out0;
assign v$G3_2816_out0 = ! v$A_4984_out0;
assign v$G3_2817_out0 = ! v$A_4985_out0;
assign v$SEL22_2923_out0 = v$A_3569_out0[8:8];
assign v$SEL13_2982_out0 = v$B_3841_out0[6:6];
assign v$SEL11_3135_out0 = v$C_4518_out0[3:3];
assign v$SEL1_3202_out0 = v$A_3569_out0[4:4];
assign v$SEL5_3239_out0 = v$A_4699_out0[5:5];
assign v$SEL9_3316_out0 = v$B_3841_out0[1:1];
assign v$SEL26_3328_out0 = v$A_4699_out0[7:7];
assign v$SEL24_3660_out0 = v$C_2732_out0[0:0];
assign v$SEL17_3824_out0 = v$A_4699_out0[0:0];
assign v$SEL11_3875_out0 = v$C_2732_out0[3:3];
assign v$SEL12_4140_out0 = v$B_3841_out0[5:5];
assign v$SEL5_4147_out0 = v$A_3569_out0[5:5];
assign v$SEL18_4246_out0 = v$B_3841_out0[3:3];
assign v$SEL9_4261_out0 = v$B_2057_out0[1:1];
assign v$11_4306_out0 = v$G6_3368_out0;
assign v$SEL21_4309_out0 = v$C_4518_out0[6:6];
assign v$SEL28_4555_out0 = v$A_3569_out0[9:9];
assign v$SEL13_4643_out0 = v$B_2057_out0[6:6];
assign v$SEL25_4720_out0 = v$C_4518_out0[2:2];
assign v$SEL7_4775_out0 = v$B_2057_out0[0:0];
assign v$SEL14_4787_out0 = v$C_2732_out0[7:7];
assign v$SEL10_4865_out0 = v$C_4518_out0[8:8];
assign v$SEL2_5056_out0 = v$A_4699_out0[6:6];
assign v$SEL14_5215_out0 = v$C_4518_out0[7:7];
assign v$G5_5361_out0 = v$A_4972_out0 && v$B_62_out0;
assign v$G5_5367_out0 = v$A_4978_out0 && v$B_68_out0;
assign v$G5_5368_out0 = v$A_4979_out0 && v$B_69_out0;
assign v$G5_5370_out0 = v$A_4981_out0 && v$B_71_out0;
assign v$G5_5373_out0 = v$A_4984_out0 && v$B_74_out0;
assign v$G5_5374_out0 = v$A_4985_out0 && v$B_75_out0;
assign v$C3_28_out0 = v$SEL11_3135_out0;
assign v$C2_198_out0 = v$SEL25_4720_out0;
assign v$A6_210_out0 = v$SEL2_604_out0;
assign v$A1_304_out0 = v$SEL16_2266_out0;
assign v$B6_346_out0 = v$SEL13_4643_out0;
assign v$A3_369_out0 = v$SEL27_918_out0;
assign v$C0_419_out0 = v$SEL24_3660_out0;
assign v$A3_491_out0 = v$SEL27_412_out0;
assign v$10_549_out0 = v$G20_319_out0;
assign v$C_640_out0 = v$G5_5361_out0;
assign v$C_646_out0 = v$G5_5367_out0;
assign v$C_647_out0 = v$G5_5368_out0;
assign v$C_649_out0 = v$G5_5370_out0;
assign v$C_652_out0 = v$G5_5373_out0;
assign v$C_653_out0 = v$G5_5374_out0;
assign v$C9_698_out0 = v$SEL30_1614_out0;
assign v$B3_705_out0 = v$SEL18_2406_out0;
assign v$G26_819_out0 = v$G22_3337_out0 && v$G23_1485_out0;
assign v$B3_877_out0 = v$SEL18_4246_out0;
assign v$A0_914_out0 = v$SEL17_993_out0;
assign v$C0_1108_out0 = v$SEL24_1408_out0;
assign v$A9_1281_out0 = v$SEL28_4555_out0;
assign v$C1_1391_out0 = v$SEL3_1663_out0;
assign v$B9_1441_out0 = v$SEL29_97_out0;
assign v$A8_1453_out0 = v$SEL22_2923_out0;
assign v$C5_1682_out0 = v$SEL4_768_out0;
assign v$C6_1683_out0 = v$SEL21_969_out0;
assign v$B1_1748_out0 = v$SEL9_4261_out0;
assign v$G21_1801_out0 = v$SEL6_1561_out0 && v$G23_1485_out0;
assign v$G0_1976_out0 = v$A_4972_out0 && v$G4_1332_out0;
assign v$G0_1982_out0 = v$A_4978_out0 && v$G4_1338_out0;
assign v$G0_1983_out0 = v$A_4979_out0 && v$G4_1339_out0;
assign v$G0_1985_out0 = v$A_4981_out0 && v$G4_1341_out0;
assign v$G0_1988_out0 = v$A_4984_out0 && v$G4_1344_out0;
assign v$G0_1989_out0 = v$A_4985_out0 && v$G4_1345_out0;
assign v$A6_2072_out0 = v$SEL2_5056_out0;
assign v$C3_2105_out0 = v$SEL11_3875_out0;
assign v$A2_2130_out0 = v$SEL15_496_out0;
assign v$A4_2221_out0 = v$SEL1_3202_out0;
assign v$B4_2250_out0 = v$SEL6_1508_out0;
assign v$C8_2449_out0 = v$SEL10_4865_out0;
assign v$B4_2468_out0 = v$SEL6_2599_out0;
assign v$G1_2519_out0 = v$G3_2804_out0 && v$B_62_out0;
assign v$G1_2525_out0 = v$G3_2810_out0 && v$B_68_out0;
assign v$G1_2526_out0 = v$G3_2811_out0 && v$B_69_out0;
assign v$G1_2528_out0 = v$G3_2813_out0 && v$B_71_out0;
assign v$G1_2531_out0 = v$G3_2816_out0 && v$B_74_out0;
assign v$G1_2532_out0 = v$G3_2817_out0 && v$B_75_out0;
assign v$B2_2646_out0 = v$SEL19_1533_out0;
assign v$B5_2656_out0 = v$SEL12_2598_out0;
assign v$B6_2663_out0 = v$SEL13_2982_out0;
assign v$A5_2706_out0 = v$SEL5_3239_out0;
assign v$A2_2729_out0 = v$SEL15_831_out0;
assign v$A4_3034_out0 = v$SEL1_1279_out0;
assign v$B8_3055_out0 = v$SEL20_1842_out0;
assign v$B1_3236_out0 = v$SEL9_3316_out0;
assign v$B7_3401_out0 = v$SEL23_9_out0;
assign v$A0_3432_out0 = v$SEL17_3824_out0;
assign v$MUX9_3446_out0 = v$11_4306_out0 ? v$C3_5358_out0 : v$MUX13_850_out0;
assign v$B2_3532_out0 = v$SEL19_1071_out0;
assign v$A1_3821_out0 = v$SEL16_1896_out0;
assign v$B7_3919_out0 = v$SEL23_585_out0;
assign v$B5_4005_out0 = v$SEL12_4140_out0;
assign v$A7_4079_out0 = v$SEL26_3328_out0;
assign v$A7_4164_out0 = v$SEL26_1764_out0;
assign v$C4_4229_out0 = v$SEL8_1504_out0;
assign v$C7_4233_out0 = v$SEL14_5215_out0;
assign v$C4_4252_out0 = v$SEL8_355_out0;
assign v$B0_4341_out0 = v$SEL7_1848_out0;
assign v$C5_4630_out0 = v$SEL4_39_out0;
assign v$A5_4739_out0 = v$SEL5_4147_out0;
assign v$C7_5135_out0 = v$SEL14_4787_out0;
assign v$_5137_out0 = { v$12_5203_out0,v$11_4306_out0 };
assign v$C6_5171_out0 = v$SEL21_4309_out0;
assign v$C2_5280_out0 = v$SEL25_1731_out0;
assign v$B0_5331_out0 = v$SEL7_4775_out0;
assign v$C1_5356_out0 = v$SEL3_1276_out0;
assign {v$A4_343_out1,v$A4_343_out0 } = v$B1_3236_out0 + v$C1_1391_out0 + v$A1_3821_out0;
assign v$G2_431_out0 = v$G0_1976_out0 || v$G1_2519_out0;
assign v$G2_437_out0 = v$G0_1982_out0 || v$G1_2525_out0;
assign v$G2_438_out0 = v$G0_1983_out0 || v$G1_2526_out0;
assign v$G2_440_out0 = v$G0_1985_out0 || v$G1_2528_out0;
assign v$G2_443_out0 = v$G0_1988_out0 || v$G1_2531_out0;
assign v$G2_444_out0 = v$G0_1989_out0 || v$G1_2532_out0;
assign {v$A4_541_out1,v$A4_541_out0 } = v$B1_1748_out0 + v$C1_5356_out0 + v$A1_304_out0;
assign {v$A1_1023_out1,v$A1_1023_out0 } = v$B4_2468_out0 + v$C4_4252_out0 + v$A4_3034_out0;
assign v$_1212_out0 = { v$C_652_out0,v$C_653_out0 };
assign {v$A1_1300_out1,v$A1_1300_out0 } = v$B4_2250_out0 + v$C4_4229_out0 + v$A4_2221_out0;
assign v$_1320_out0 = { v$C6_3912_out0,v$C_647_out0 };
assign v$_1323_out0 = { v$C7_825_out0,v$C_646_out0 };
assign {v$A9_1329_out1,v$A9_1329_out0 } = v$B5_2656_out0 + v$C5_1682_out0 + v$A5_2706_out0;
assign {v$A8_1629_out1,v$A8_1629_out0 } = v$B8_3055_out0 + v$C8_2449_out0 + v$A8_1453_out0;
assign {v$A6_1657_out1,v$A6_1657_out0 } = v$B6_2663_out0 + v$C6_5171_out0 + v$A6_210_out0;
assign {v$A5_1759_out1,v$A5_1759_out0 } = v$B2_3532_out0 + v$C2_5280_out0 + v$A2_2130_out0;
assign v$9_2616_out0 = v$G21_1801_out0;
assign v$G24_2701_out0 = v$SEL7_1406_out0 && v$G26_819_out0;
assign v$G42_2708_out0 = v$G40_2290_out0 && v$G26_819_out0;
assign {v$A2_3190_out1,v$A2_3190_out0 } = v$B3_705_out0 + v$C3_2105_out0 + v$A3_491_out0;
assign {v$A10_3266_out1,v$A10_3266_out0 } = v$B9_1441_out0 + v$C9_698_out0 + v$A9_1281_out0;
assign {v$A7_3669_out1,v$A7_3669_out0 } = v$B0_4341_out0 + v$C0_1108_out0 + v$A0_914_out0;
assign {v$A3_3731_out1,v$A3_3731_out0 } = v$B7_3401_out0 + v$C7_5135_out0 + v$A7_4079_out0;
assign {v$A9_3764_out1,v$A9_3764_out0 } = v$B5_4005_out0 + v$C5_4630_out0 + v$A5_4739_out0;
assign {v$A7_3868_out1,v$A7_3868_out0 } = v$B0_5331_out0 + v$C0_419_out0 + v$A0_3432_out0;
assign v$MUX12_3906_out0 = v$10_549_out0 ? v$C4_1032_out0 : v$MUX9_3446_out0;
assign {v$A6_4050_out1,v$A6_4050_out0 } = v$B6_346_out0 + v$C6_1683_out0 + v$A6_2072_out0;
assign {v$A2_4329_out1,v$A2_4329_out0 } = v$B3_877_out0 + v$C3_28_out0 + v$A3_369_out0;
assign {v$A5_4640_out1,v$A5_4640_out0 } = v$B2_2646_out0 + v$C2_198_out0 + v$A2_2729_out0;
assign {v$A3_5327_out1,v$A3_5327_out0 } = v$B7_3919_out0 + v$C7_4233_out0 + v$A7_4164_out0;
assign v$S12_101_out0 = v$A5_4640_out1;
assign v$S15_542_out0 = v$A9_1329_out1;
assign v$S19_569_out0 = v$A10_3266_out1;
assign v$MUX10_590_out0 = v$9_2616_out0 ? v$C5_4465_out0 : v$MUX12_3906_out0;
assign v$S14_668_out0 = v$A1_1300_out1;
assign v$S14_753_out0 = v$A1_1023_out1;
assign v$_776_out0 = { v$_1212_out0,v$C_640_out0 };
assign v$S13_852_out0 = v$A2_4329_out1;
assign v$S07_887_out0 = v$A3_5327_out0;
assign v$S10_939_out0 = v$A7_3669_out1;
assign v$S01_1062_out0 = v$A4_343_out0;
assign v$_1070_out0 = { v$10_549_out0,v$9_2616_out0 };
assign v$S13_1157_out0 = v$A2_3190_out1;
assign v$S02_1187_out0 = v$A5_1759_out0;
assign v$G41_1468_out0 = v$G45_2793_out0 && v$G42_2708_out0;
assign v$S08_1590_out0 = v$A8_1629_out0;
assign v$S09_1937_out0 = v$A10_3266_out0;
assign v$8_1973_out0 = v$G24_2701_out0;
assign v$S04_2279_out0 = v$A1_1300_out0;
assign v$G43_2435_out0 = v$SEL14_1155_out0 && v$G42_2708_out0;
assign v$S18_2437_out0 = v$A8_1629_out1;
assign v$S03_2845_out0 = v$A2_4329_out0;
assign v$S00_2884_out0 = v$A7_3868_out0;
assign v$S06_3112_out0 = v$A6_1657_out0;
assign v$S11_3141_out0 = v$A4_343_out1;
assign v$S15_3217_out0 = v$A9_3764_out1;
assign v$S16_3242_out0 = v$A6_4050_out1;
assign v$S10_3263_out0 = v$A7_3868_out1;
assign v$S06_3373_out0 = v$A6_4050_out0;
assign v$S02_3391_out0 = v$A5_4640_out0;
assign v$S05_3458_out0 = v$A9_1329_out0;
assign v$S11_3803_out0 = v$A4_541_out1;
assign v$S03_4045_out0 = v$A2_3190_out0;
assign v$S17_4091_out0 = v$A3_5327_out1;
assign v$S17_4121_out0 = v$A3_3731_out1;
assign v$S_4177_out0 = v$G2_431_out0;
assign v$S_4183_out0 = v$G2_437_out0;
assign v$S_4184_out0 = v$G2_438_out0;
assign v$S_4186_out0 = v$G2_440_out0;
assign v$S_4189_out0 = v$G2_443_out0;
assign v$S_4190_out0 = v$G2_444_out0;
assign v$S00_4440_out0 = v$A7_3669_out0;
assign v$S12_4495_out0 = v$A5_1759_out1;
assign v$S16_4695_out0 = v$A6_1657_out1;
assign v$S04_4731_out0 = v$A1_1023_out0;
assign v$S05_4887_out0 = v$A9_3764_out0;
assign v$S07_5042_out0 = v$A3_3731_out0;
assign v$S01_5221_out0 = v$A4_541_out0;
assign v$_175_out0 = { v$S08_1590_out0,v$S09_1937_out0 };
assign v$_237_out0 = { v$S18_2437_out0,v$S19_569_out0 };
assign v$_404_out0 = { v$S16_3242_out0,v$S17_4121_out0 };
assign v$_717_out0 = { v$S10_3263_out0,v$S11_3803_out0 };
assign v$_944_out0 = { v$S02_3391_out0,v$S03_2845_out0 };
assign v$_1164_out0 = { v$S00_4440_out0,v$S01_1062_out0 };
assign v$_1593_out0 = { v$SEL48_4857_out0,v$S_4184_out0 };
assign v$_1723_out0 = { v$S06_3373_out0,v$S07_5042_out0 };
assign v$_1878_out0 = { v$S04_4731_out0,v$S05_3458_out0 };
assign v$MUX11_1882_out0 = v$8_1973_out0 ? v$C6_4824_out0 : v$MUX10_590_out0;
assign v$_1889_out0 = { v$S16_4695_out0,v$S17_4091_out0 };
assign v$_2402_out0 = { v$S00_2884_out0,v$S01_5221_out0 };
assign v$_2630_out0 = { v$S_4189_out0,v$S_4190_out0 };
assign v$G48_2727_out0 = v$G46_561_out0 && v$G41_1468_out0;
assign v$_2735_out0 = { v$S10_939_out0,v$S11_3141_out0 };
assign v$_3108_out0 = { v$S14_668_out0,v$S15_3217_out0 };
assign v$G44_3211_out0 = v$SEL13_3457_out0 && v$G41_1468_out0;
assign v$_3576_out0 = { v$S06_3112_out0,v$S07_887_out0 };
assign v$_3600_out0 = { v$_5137_out0,v$_1070_out0 };
assign v$_3815_out0 = { v$S12_101_out0,v$S13_852_out0 };
assign v$_4438_out0 = { v$S14_753_out0,v$S15_542_out0 };
assign v$_4491_out0 = { v$S02_1187_out0,v$S03_4045_out0 };
assign v$_4769_out0 = { v$S12_4495_out0,v$S13_1157_out0 };
assign v$_4863_out0 = { v$_5278_out0,v$S_4183_out0 };
assign v$_4879_out0 = { v$S04_2279_out0,v$S05_4887_out0 };
assign v$7_4953_out0 = v$G43_2435_out0;
assign v$_376_out0 = { v$_4438_out0,v$_404_out0 };
assign v$_532_out0 = { v$_2630_out0,v$S_4177_out0 };
assign v$_1421_out0 = { v$_2735_out0,v$_3815_out0 };
assign v$_1671_out0 = { v$_4879_out0,v$_3576_out0 };
assign v$_1747_out0 = { v$8_1973_out0,v$7_4953_out0 };
assign v$_2018_out0 = { v$_3108_out0,v$_1889_out0 };
assign v$_2074_out0 = { v$_1164_out0,v$_944_out0 };
assign v$_2192_out0 = { v$_717_out0,v$_4769_out0 };
assign v$MUX8_2409_out0 = v$7_4953_out0 ? v$C7_1909_out0 : v$MUX11_1882_out0;
assign v$_2705_out0 = { v$_2402_out0,v$_4491_out0 };
assign v$G49_3414_out0 = v$SEL16_4040_out0 && v$G48_2727_out0;
assign v$6_3497_out0 = v$G44_3211_out0;
assign v$_3725_out0 = { v$_1878_out0,v$_1723_out0 };
assign v$G47_4375_out0 = v$G51_3597_out0 && v$G48_2727_out0;
assign v$G50_248_out0 = v$SEL15_469_out0 && v$G47_4375_out0;
assign v$_688_out0 = { v$_1671_out0,v$_175_out0 };
assign v$G54_2010_out0 = v$G52_303_out0 && v$G47_4375_out0;
assign v$MUX6_3119_out0 = v$6_3497_out0 ? v$C8_2635_out0 : v$MUX8_2409_out0;
assign v$_3435_out0 = { v$_2705_out0,v$_3725_out0 };
assign v$_3537_out0 = { v$_2192_out0,v$_376_out0 };
assign v$_4057_out0 = { v$_2018_out0,v$_237_out0 };
assign v$5_4221_out0 = v$G49_3414_out0;
assign v$4_1202_out0 = v$G50_248_out0;
assign v$MUX5_1752_out0 = v$5_4221_out0 ? v$C9_2797_out0 : v$MUX6_3119_out0;
assign v$S2_2248_out0 = v$_3537_out0;
assign v$G53_2297_out0 = v$G57_4885_out0 && v$G54_2010_out0;
assign v$S1_2964_out0 = v$_3435_out0;
assign v$_3039_out0 = { v$_1421_out0,v$_4057_out0 };
assign v$G55_3409_out0 = v$SEL18_26_out0 && v$G54_2010_out0;
assign v$_3609_out0 = { v$_2074_out0,v$_688_out0 };
assign v$_4790_out0 = { v$6_3497_out0,v$5_4221_out0 };
assign v$_1_out0 = { v$S_4186_out0,v$S1_2964_out0 };
assign v$MUX7_526_out0 = v$4_1202_out0 ? v$C10_1969_out0 : v$MUX5_1752_out0;
assign v$G56_2856_out0 = v$SEL17_3946_out0 && v$G53_2297_out0;
assign v$_3122_out0 = { v$_1747_out0,v$_4790_out0 };
assign v$S1_4206_out0 = v$_3609_out0;
assign v$S2_4316_out0 = v$_3039_out0;
assign v$_4320_out0 = { v$C_649_out0,v$S2_2248_out0 };
assign v$3_4628_out0 = v$G55_3409_out0;
assign v$G60_5428_out0 = v$G58_4585_out0 && v$G53_2297_out0;
assign v$_22_out0 = { v$4_1202_out0,v$3_4628_out0 };
assign v$MUX4_726_out0 = v$3_4628_out0 ? v$C11_3343_out0 : v$MUX7_526_out0;
assign v$G63_823_out0 = v$G62_4943_out0 && v$G60_5428_out0;
assign v$_2316_out0 = { v$_3600_out0,v$_3122_out0 };
assign v$_2578_out0 = { v$_4863_out0,v$_1_out0 };
assign v$2_2919_out0 = v$G56_2856_out0;
assign v$_3442_out0 = { v$_1320_out0,v$S2_4316_out0 };
assign v$_3813_out0 = { v$_1323_out0,v$_4320_out0 };
assign v$G61_3943_out0 = v$SEL20_2272_out0 && v$G60_5428_out0;
assign v$_4940_out0 = { v$S1_4206_out0,v$SEL90_2866_out0 };
assign v$_19_out0 = { v$_3442_out0,v$SEL47_4498_out0 };
assign v$G65_131_out0 = v$G66_558_out0 && v$G63_823_out0;
assign v$_1370_out0 = { v$_3813_out0,v$_776_out0 };
assign v$_1716_out0 = { v$_2578_out0,v$_532_out0 };
assign v$G64_2690_out0 = v$G63_823_out0 && v$SEL21_2093_out0;
assign v$MUX3_2998_out0 = v$2_2919_out0 ? v$C12_2311_out0 : v$MUX4_726_out0;
assign v$1_3429_out0 = v$G61_3943_out0;
assign v$_5179_out0 = { v$_1593_out0,v$_4940_out0 };
assign v$_363_out0 = { v$2_2919_out0,v$1_3429_out0 };
assign v$M0_573_out0 = v$_5179_out0;
assign v$M1_973_out0 = v$_19_out0;
assign v$MUX2_1040_out0 = v$1_3429_out0 ? v$C13_1293_out0 : v$MUX3_2998_out0;
assign v$M2_1829_out0 = v$_1716_out0;
assign v$M3_3543_out0 = v$_1370_out0;
assign v$0_4365_out0 = v$G64_2690_out0;
assign v$SERIESCONNECT_4606_out0 = v$G65_131_out0;
assign v$SEL75_158_out0 = v$M0_573_out0[13:5];
assign v$SEL72_215_out0 = v$M2_1829_out0[15:15];
assign v$SEL87_244_out0 = v$M3_3543_out0[9:9];
assign v$_485_out0 = { v$0_4365_out0,v$1_3429_out0 };
assign v$SEL67_815_out0 = v$M1_973_out0[3:3];
assign v$SEL69_824_out0 = v$M2_1829_out0[13:5];
assign v$_1003_out0 = { v$_22_out0,v$_363_out0 };
assign v$SEL89_1033_out0 = v$M3_3543_out0[8:7];
assign v$SEL74_1540_out0 = v$M0_573_out0[4:4];
assign v$SEL80_1577_out0 = v$M1_973_out0[14:14];
assign v$SEL77_2323_out0 = v$M1_973_out0[15:15];
assign v$SEL83_2369_out0 = v$M3_3543_out0[19:10];
assign v$SEL70_2638_out0 = v$M1_973_out0[4:4];
assign v$SEL82_2669_out0 = v$M2_1829_out0[16:16];
assign v$MUX1_2933_out0 = v$0_4365_out0 ? v$C14_2741_out0 : v$MUX2_1040_out0;
assign v$SEL71_3374_out0 = v$M2_1829_out0[14:14];
assign v$SEL68_3726_out0 = v$M0_573_out0[2:0];
assign v$SEL81_3767_out0 = v$M2_1829_out0[18:17];
assign v$SEL78_4371_out0 = v$M0_573_out0[3:3];
assign v$SEL73_4687_out0 = v$M1_973_out0[13:5];
assign v$X1_4916_out0 = v$SERIESCONNECT_4606_out0;
assign v$B_64_out0 = v$SEL80_1577_out0;
assign v$B_65_out0 = v$SEL77_2323_out0;
assign v$B_70_out0 = v$SEL67_815_out0;
assign v$B_76_out0 = v$SEL70_2638_out0;
assign v$SHIFTNUMBER_337_out0 = v$MUX1_2933_out0;
assign v$_1180_out0 = { v$_485_out0,v$2_2919_out0 };
assign v$_2254_out0 = { v$C13_274_out0,v$SEL89_1033_out0 };
assign v$C_3601_out0 = v$SEL75_158_out0;
assign v$_3607_out0 = { v$_1003_out0,v$0_4365_out0 };
assign v$A_3704_out0 = v$SEL69_824_out0;
assign v$B_3711_out0 = v$SEL73_4687_out0;
assign v$B_3842_out0 = v$SEL83_2369_out0;
assign v$A_4973_out0 = v$SEL87_244_out0;
assign v$A_4974_out0 = v$SEL71_3374_out0;
assign v$A_4975_out0 = v$SEL72_215_out0;
assign v$A_4980_out0 = v$SEL78_4371_out0;
assign v$A_4986_out0 = v$SEL74_1540_out0;
assign v$SEL29_98_out0 = v$B_3842_out0[9:9];
assign v$SEL3_357_out0 = v$A_3704_out0[4:4];
assign v$SEL23_586_out0 = v$B_3842_out0[7:7];
assign v$SEL2_739_out0 = v$A_3704_out0[6:6];
assign v$SEL21_754_out0 = v$C_3601_out0[1:1];
assign v$SEL22_958_out0 = v$C_3601_out0[5:5];
assign v$SEL6_1041_out0 = v$A_3704_out0[5:5];
assign v$SEL10_1158_out0 = v$B_3711_out0[4:4];
assign v$G4_1334_out0 = ! v$B_64_out0;
assign v$G4_1335_out0 = ! v$B_65_out0;
assign v$G4_1340_out0 = ! v$B_70_out0;
assign v$G4_1346_out0 = ! v$B_76_out0;
assign v$SEL15_1363_out0 = v$B_3711_out0[0:0];
assign v$SEL19_1486_out0 = v$C_3601_out0[4:4];
assign v$SEL14_1491_out0 = v$B_3711_out0[1:1];
assign v$SEL6_1509_out0 = v$B_3842_out0[4:4];
assign v$SEL19_1534_out0 = v$B_3842_out0[2:2];
assign v$SEL26_1706_out0 = v$C_3601_out0[8:8];
assign v$SEL24_1791_out0 = v$C_3601_out0[3:3];
assign v$SEL20_1843_out0 = v$B_3842_out0[8:8];
assign v$SEL7_1849_out0 = v$B_3842_out0[0:0];
assign v$G0_1977_out0 = v$A_4973_out0 && v$G4_1333_out0;
assign v$SEL12_2081_out0 = v$B_3711_out0[5:5];
assign v$_2425_out0 = { v$_2316_out0,v$_3607_out0 };
assign v$SEL11_2549_out0 = v$B_3711_out0[6:6];
assign v$SEL27_2607_out0 = v$C_3601_out0[7:7];
assign v$G3_2805_out0 = ! v$A_4973_out0;
assign v$G3_2806_out0 = ! v$A_4974_out0;
assign v$G3_2807_out0 = ! v$A_4975_out0;
assign v$G3_2812_out0 = ! v$A_4980_out0;
assign v$G3_2818_out0 = ! v$A_4986_out0;
assign v$SEL13_2983_out0 = v$B_3842_out0[6:6];
assign v$SEL4_3161_out0 = v$A_3704_out0[2:2];
assign v$SEL1_3305_out0 = v$A_3704_out0[1:1];
assign v$SEL9_3317_out0 = v$B_3842_out0[1:1];
assign v$SEL9_3386_out0 = v$A_3704_out0[0:0];
assign v$SEL18_3449_out0 = v$B_3711_out0[3:3];
assign v$_3623_out0 = { v$_1180_out0,v$3_4628_out0 };
assign v$SEL13_3869_out0 = v$B_3711_out0[2:2];
assign v$SEL16_3937_out0 = v$B_3711_out0[8:8];
assign v$SEL23_3968_out0 = v$C_3601_out0[6:6];
assign v$SEL5_4029_out0 = v$A_3704_out0[8:8];
assign v$SEL12_4141_out0 = v$B_3842_out0[5:5];
assign v$SEL18_4247_out0 = v$B_3842_out0[3:3];
assign v$SEL17_4471_out0 = v$B_3711_out0[7:7];
assign v$SEL20_4543_out0 = v$C_3601_out0[0:0];
assign v$SEL25_4655_out0 = v$C_3601_out0[2:2];
assign v$SEL8_4725_out0 = v$A_3704_out0[7:7];
assign v$SHIFTNUMBER_5177_out0 = v$SHIFTNUMBER_337_out0;
assign v$SEL7_5191_out0 = v$A_3704_out0[3:3];
assign v$G5_5362_out0 = v$A_4973_out0 && v$B_63_out0;
assign v$G5_5363_out0 = v$A_4974_out0 && v$B_64_out0;
assign v$G5_5364_out0 = v$A_4975_out0 && v$B_65_out0;
assign v$G5_5369_out0 = v$A_4980_out0 && v$B_70_out0;
assign v$G5_5375_out0 = v$A_4986_out0 && v$B_76_out0;
assign v$A5_50_out0 = v$SEL6_1041_out0;
assign v$A2_312_out0 = v$SEL4_3161_out0;
assign v$A0_550_out0 = v$SEL9_3386_out0;
assign v$C_641_out0 = v$G5_5362_out0;
assign v$C_642_out0 = v$G5_5363_out0;
assign v$C_643_out0 = v$G5_5364_out0;
assign v$C_648_out0 = v$G5_5369_out0;
assign v$C_654_out0 = v$G5_5375_out0;
assign v$A1_731_out0 = v$SEL1_3305_out0;
assign v$B2_764_out0 = v$SEL13_3869_out0;
assign v$B3_878_out0 = v$SEL18_4247_out0;
assign v$A3_1052_out0 = v$SEL7_5191_out0;
assign v$B9_1442_out0 = v$SEL29_98_out0;
assign v$A8_1556_out0 = v$SEL5_4029_out0;
assign v$B4_1867_out0 = v$SEL10_1158_out0;
assign v$G0_1978_out0 = v$A_4974_out0 && v$G4_1334_out0;
assign v$G0_1979_out0 = v$A_4975_out0 && v$G4_1335_out0;
assign v$G0_1984_out0 = v$A_4980_out0 && v$G4_1340_out0;
assign v$G0_1990_out0 = v$A_4986_out0 && v$G4_1346_out0;
assign v$B7_2160_out0 = v$SEL17_4471_out0;
assign v$B8_2201_out0 = v$SEL16_3937_out0;
assign v$B4_2251_out0 = v$SEL6_1509_out0;
assign v$C7_2317_out0 = v$SEL27_2607_out0;
assign v$A4_2442_out0 = v$SEL3_357_out0;
assign v$G1_2520_out0 = v$G3_2805_out0 && v$B_63_out0;
assign v$G1_2521_out0 = v$G3_2806_out0 && v$B_64_out0;
assign v$G1_2522_out0 = v$G3_2807_out0 && v$B_65_out0;
assign v$G1_2527_out0 = v$G3_2812_out0 && v$B_70_out0;
assign v$G1_2533_out0 = v$G3_2818_out0 && v$B_76_out0;
assign v$B2_2647_out0 = v$SEL19_1534_out0;
assign v$B6_2664_out0 = v$SEL13_2983_out0;
assign v$C6_2674_out0 = v$SEL23_3968_out0;
assign v$B5_3027_out0 = v$SEL12_2081_out0;
assign v$B8_3056_out0 = v$SEL20_1843_out0;
assign v$_3087_out0 = { v$SHIFTNUMBER_5177_out0,v$C18_1516_out0 };
assign v$B1_3237_out0 = v$SEL9_3317_out0;
assign v$C4_3418_out0 = v$SEL19_1486_out0;
assign v$C5_3631_out0 = v$SEL22_958_out0;
assign v$C1_3691_out0 = v$SEL21_754_out0;
assign v$A6_3768_out0 = v$SEL2_739_out0;
assign v$B7_3920_out0 = v$SEL23_586_out0;
assign v$C2_3989_out0 = v$SEL25_4655_out0;
assign v$B5_4006_out0 = v$SEL12_4141_out0;
assign v$B0_4342_out0 = v$SEL7_1849_out0;
assign v$_4451_out0 = { v$_3623_out0,v$4_1202_out0 };
assign v$A7_4559_out0 = v$SEL8_4725_out0;
assign v$_4653_out0 = { v$SHIFTNUMBER_5177_out0,v$C21_4967_out0 };
assign v$C3_4732_out0 = v$SEL24_1791_out0;
assign v$B6_4850_out0 = v$SEL11_2549_out0;
assign v$C8_4923_out0 = v$SEL26_1706_out0;
assign v$B3_5122_out0 = v$SEL18_3449_out0;
assign v$OUTPUTSHIFT_5151_out0 = v$_2425_out0;
assign v$B0_5313_out0 = v$SEL15_1363_out0;
assign v$B1_5322_out0 = v$SEL14_1491_out0;
assign v$C0_5419_out0 = v$SEL20_4543_out0;
assign {v$A4_344_out1,v$A4_344_out0 } = v$B1_3237_out0 + v$C1_1392_out0 + v$A1_3822_out0;
assign v$G2_432_out0 = v$G0_1977_out0 || v$G1_2520_out0;
assign v$G2_433_out0 = v$G0_1978_out0 || v$G1_2521_out0;
assign v$G2_434_out0 = v$G0_1979_out0 || v$G1_2522_out0;
assign v$G2_439_out0 = v$G0_1984_out0 || v$G1_2527_out0;
assign v$G2_445_out0 = v$G0_1990_out0 || v$G1_2533_out0;
assign {v$A4_519_out1,v$A4_519_out0 } = v$B4_1867_out0 + v$C4_3418_out0 + v$A4_2442_out0;
assign v$OUTPUTSHIFT_1089_out0 = v$OUTPUTSHIFT_5151_out0;
assign {v$A6_1090_out1,v$A6_1090_out0 } = v$B3_5122_out0 + v$C3_4732_out0 + v$A3_1052_out0;
assign v$_1211_out0 = { v$_4451_out0,v$5_4221_out0 };
assign {v$A1_1301_out1,v$A1_1301_out0 } = v$B4_2251_out0 + v$C4_4230_out0 + v$A4_2222_out0;
assign {v$A8_1630_out1,v$A8_1630_out0 } = v$B8_3056_out0 + v$C8_2450_out0 + v$A8_1454_out0;
assign {v$A6_1658_out1,v$A6_1658_out0 } = v$B6_2664_out0 + v$C6_5172_out0 + v$A6_211_out0;
assign {v$A7_1862_out1,v$A7_1862_out0 } = v$B7_2160_out0 + v$C7_2317_out0 + v$A7_4559_out0;
assign {v$A2_2602_out1,v$A2_2602_out0 } = v$B1_5322_out0 + v$C1_3691_out0 + v$A1_731_out0;
assign {v$A3_2871_out1,v$A3_2871_out0 } = v$B2_764_out0 + v$C2_3989_out0 + v$A2_312_out0;
assign v$_2926_out0 = { v$C_643_out0,v$SEL81_3767_out0 };
assign v$_2944_out0 = { v$C12_45_out0,v$C_641_out0 };
assign {v$A10_3267_out1,v$A10_3267_out0 } = v$B9_1442_out0 + v$C9_699_out0 + v$A9_1282_out0;
assign v$XOR1_3486_out0 = v$_3087_out0 ^ v$C15_3897_out0;
assign v$SHIFTNUMBER5_3520_out0 = v$_4653_out0;
assign {v$A7_3670_out1,v$A7_3670_out0 } = v$B0_4342_out0 + v$C0_1109_out0 + v$A0_915_out0;
assign {v$A8_3700_out1,v$A8_3700_out0 } = v$B6_4850_out0 + v$C6_2674_out0 + v$A6_3768_out0;
assign {v$A1_3715_out1,v$A1_3715_out0 } = v$B0_5313_out0 + v$C0_5419_out0 + v$A0_550_out0;
assign {v$A9_3765_out1,v$A9_3765_out0 } = v$B5_4006_out0 + v$C5_4631_out0 + v$A5_4740_out0;
assign {v$A2_4330_out1,v$A2_4330_out0 } = v$B3_878_out0 + v$C3_29_out0 + v$A3_370_out0;
assign {v$A9_4399_out1,v$A9_4399_out0 } = v$B8_2201_out0 + v$C8_4923_out0 + v$A8_1556_out0;
assign v$_4542_out0 = { v$C11_3383_out0,v$C_648_out0 };
assign {v$A5_4641_out1,v$A5_4641_out0 } = v$B2_2647_out0 + v$C2_199_out0 + v$A2_2730_out0;
assign {v$A5_5011_out1,v$A5_5011_out0 } = v$B5_3027_out0 + v$C5_3631_out0 + v$A5_50_out0;
assign {v$A3_5328_out1,v$A3_5328_out0 } = v$B7_3920_out0 + v$C7_4234_out0 + v$A7_4165_out0;
assign v$S12_102_out0 = v$A5_4641_out1;
assign v$_161_out0 = { v$_1211_out0,v$6_3497_out0 };
assign v$S01_191_out0 = v$A2_2602_out0;
assign v$S15_458_out0 = v$A5_5011_out1;
assign v$S19_570_out0 = v$A10_3267_out1;
assign v$S14_669_out0 = v$A1_1301_out1;
assign v$S13_853_out0 = v$A2_4330_out1;
assign v$S07_888_out0 = v$A3_5328_out0;
assign v$S04_927_out0 = v$A4_519_out0;
assign v$S10_940_out0 = v$A7_3670_out1;
assign v$S01_1063_out0 = v$A4_344_out0;
assign v$S02_1072_out0 = v$A3_2871_out0;
assign v$S00_1128_out0 = v$A1_3715_out0;
assign v$S07_1254_out0 = v$A7_1862_out0;
assign v$S08_1591_out0 = v$A8_1630_out0;
assign v$S09_1938_out0 = v$A10_3267_out0;
assign v$S18_1961_out0 = v$A9_4399_out1;
assign {v$A1_2126_out1,v$A1_2126_out0 } = v$_2024_out0 + v$XOR1_3486_out0 + v$C14_4933_out0;
assign v$S04_2280_out0 = v$A1_1301_out0;
assign v$S18_2438_out0 = v$A8_1630_out1;
assign v$S11_2561_out0 = v$A2_2602_out1;
assign v$S03_2846_out0 = v$A2_4330_out0;
assign v$S17_2861_out0 = v$A7_1862_out1;
assign v$S05_2988_out0 = v$A5_5011_out0;
assign v$S03_3014_out0 = v$A6_1090_out0;
assign v$S06_3113_out0 = v$A6_1658_out0;
assign v$S11_3142_out0 = v$A4_344_out1;
assign v$S15_3218_out0 = v$A9_3765_out1;
assign v$S14_3379_out0 = v$A4_519_out1;
assign v$S02_3392_out0 = v$A5_4641_out0;
assign v$S13_3436_out0 = v$A6_1090_out1;
assign v$S10_3471_out0 = v$A1_3715_out1;
assign v$S17_4092_out0 = v$A3_5328_out1;
assign v$S_4178_out0 = v$G2_432_out0;
assign v$S_4179_out0 = v$G2_433_out0;
assign v$S_4180_out0 = v$G2_434_out0;
assign v$S_4185_out0 = v$G2_439_out0;
assign v$S_4191_out0 = v$G2_445_out0;
assign v$S06_4367_out0 = v$A8_3700_out0;
assign v$_4393_out0 = { v$C_642_out0,v$_2926_out0 };
assign v$S00_4441_out0 = v$A7_3670_out0;
assign v$S16_4696_out0 = v$A6_1658_out1;
assign v$S12_4798_out0 = v$A3_2871_out1;
assign v$S05_4888_out0 = v$A9_3765_out0;
assign v$S16_4891_out0 = v$A8_3700_out1;
assign v$S08_5271_out0 = v$A9_4399_out0;
assign v$_176_out0 = { v$S08_1591_out0,v$S09_1938_out0 };
assign v$_238_out0 = { v$S18_2438_out0,v$S19_570_out0 };
assign v$_839_out0 = { v$S10_3471_out0,v$S11_2561_out0 };
assign v$_863_out0 = v$A1_2126_out0[4:0];
assign v$_863_out1 = v$A1_2126_out0[5:1];
assign v$_945_out0 = { v$S02_3392_out0,v$S03_2846_out0 };
assign v$COUT_1151_out0 = v$A1_2126_out1;
assign v$_1165_out0 = { v$S00_4441_out0,v$S01_1063_out0 };
assign v$_1430_out0 = { v$S04_927_out0,v$S05_2988_out0 };
assign v$_1607_out0 = { v$S02_1072_out0,v$S03_3014_out0 };
assign v$_1890_out0 = { v$S16_4696_out0,v$S17_4092_out0 };
assign v$_2353_out0 = { v$S12_4798_out0,v$S13_3436_out0 };
assign v$EQ15_2421_out0 = v$A1_2126_out0 == 6'h0;
assign v$_2736_out0 = { v$S10_940_out0,v$S11_3142_out0 };
assign v$_2977_out0 = { v$S16_4891_out0,v$S17_2861_out0 };
assign v$_3109_out0 = { v$S14_669_out0,v$S15_3218_out0 };
assign v$_3360_out0 = { v$_161_out0,v$7_4953_out0 };
assign v$_3577_out0 = { v$S06_3113_out0,v$S07_888_out0 };
assign v$_3586_out0 = { v$S_4180_out0,v$SEL82_2669_out0 };
assign v$_3590_out0 = { v$_2254_out0,v$S_4178_out0 };
assign v$_3624_out0 = { v$S06_4367_out0,v$S07_1254_out0 };
assign v$_3637_out0 = { v$S00_1128_out0,v$S01_191_out0 };
assign v$_3816_out0 = { v$S12_102_out0,v$S13_853_out0 };
assign v$_4126_out0 = { v$S14_3379_out0,v$S15_458_out0 };
assign v$_4717_out0 = { v$SEL68_3726_out0,v$S_4185_out0 };
assign v$_4880_out0 = { v$S04_2280_out0,v$S05_4888_out0 };
assign v$_107_out0 = { v$_3360_out0,v$8_1973_out0 };
assign v$EQ16_330_out0 = v$_863_out1 == 1'h0;
assign {v$A2_528_out1,v$A2_528_out0 } = v$_863_out0 + v$C20_4877_out0 + v$DETECT1_1926_out0;
assign v$_1419_out0 = { v$S_4179_out0,v$_3586_out0 };
assign v$_1422_out0 = { v$_2736_out0,v$_3816_out0 };
assign v$_1603_out0 = { v$_4126_out0,v$_2977_out0 };
assign v$_1672_out0 = { v$_4880_out0,v$_3577_out0 };
assign v$_2019_out0 = { v$_3109_out0,v$_1890_out0 };
assign v$_2075_out0 = { v$_1165_out0,v$_945_out0 };
assign v$_2658_out0 = { v$_1430_out0,v$_3624_out0 };
assign v$_4157_out0 = { v$_3637_out0,v$_1607_out0 };
assign v$_4753_out0 = { v$_839_out0,v$_2353_out0 };
assign v$EQUAL_5339_out0 = v$EQ15_2421_out0;
assign v$DIFFERENCE_133_out0 = v$A2_528_out0;
assign v$_689_out0 = { v$_1672_out0,v$_176_out0 };
assign v$_1291_out0 = { v$_107_out0,v$9_2616_out0 };
assign v$_2462_out0 = { v$_2658_out0,v$S08_5271_out0 };
assign v$EXPOBIGGER_2483_out0 = v$EQ16_330_out0;
assign v$NOTUSE_3678_out0 = v$A2_528_out1;
assign v$_4058_out0 = { v$_2019_out0,v$_238_out0 };
assign v$_4322_out0 = { v$_1603_out0,v$S18_1961_out0 };
assign v$MUX14_142_out0 = v$EXPOBIGGER_2483_out0 ? v$SHIFTNUMBER5_3520_out0 : v$MUX23_5205_out0;
assign v$_216_out0 = { v$_4753_out0,v$_4322_out0 };
assign v$MUX16_908_out0 = v$EQUAL_5339_out0 ? v$MUX22_3031_out0 : v$DIFFERENCE_133_out0;
assign v$_934_out0 = { v$_1291_out0,v$10_549_out0 };
assign v$_3040_out0 = { v$_1422_out0,v$_4058_out0 };
assign v$_3610_out0 = { v$_2075_out0,v$_689_out0 };
assign v$_3864_out0 = { v$_4157_out0,v$_2462_out0 };
assign v$SHIFTNUMBER_672_out0 = v$MUX14_142_out0;
assign v$S0_1259_out0 = v$_3864_out0;
assign v$S1_4207_out0 = v$_3610_out0;
assign v$S1_4224_out0 = v$_216_out0;
assign v$S2_4317_out0 = v$_3040_out0;
assign v$MUX15_5223_out0 = v$EXPOBIGGER_2483_out0 ? v$MUX16_908_out0 : v$C16_206_out0;
assign v$_5399_out0 = { v$_934_out0,v$11_4306_out0 };
assign v$_10_out0 = { v$_2944_out0,v$S2_4317_out0 };
assign v$_601_out0 = { v$_5399_out0,v$12_5203_out0 };
assign v$SHIFTNUMBER1_611_out0 = v$SHIFTNUMBER_672_out0;
assign v$SEL3_1482_out0 = v$SHIFTNUMBER_672_out0[3:3];
assign v$SEL5_1596_out0 = v$SHIFTNUMBER_672_out0[2:2];
assign v$NEWEXPONENT_1711_out0 = v$MUX15_5223_out0;
assign v$SEL4_3355_out0 = v$SHIFTNUMBER_672_out0[4:4];
assign v$_3916_out0 = { v$S_4191_out0,v$S0_1259_out0 };
assign v$_4443_out0 = { v$C_654_out0,v$S1_4224_out0 };
assign v$SEL1_4771_out0 = v$SHIFTNUMBER_672_out0[0:0];
assign v$SEL2_4934_out0 = v$SHIFTNUMBER_672_out0[1:1];
assign v$_5251_out0 = { v$S1_4207_out0,v$SEL88_4558_out0 };
assign v$_1099_out0 = { v$_3590_out0,v$_5251_out0 };
assign v$OUTPUT_1821_out0 = v$_601_out0;
assign v$MUX20_3019_out0 = v$SEL4_3355_out0 ? v$C25_3774_out0 : v$INPUT_3065_out0;
assign v$_3020_out0 = { v$_4542_out0,v$_4443_out0 };
assign v$N3_3326_out0 = v$_10_out0;
assign v$_4072_out0 = { v$_4717_out0,v$_3916_out0 };
assign v$NEWEXPO_4492_out0 = v$NEWEXPONENT_1711_out0;
assign v$SHIFTNUM_5219_out0 = v$SHIFTNUMBER1_611_out0;
assign v$_500_out0 = { v$_3020_out0,v$_4393_out0 };
assign v$_735_out0 = { v$_4072_out0,v$_1419_out0 };
assign v$N2_820_out0 = v$_1099_out0;
assign v$X_1476_out0 = v$OUTPUT_1821_out0;
assign v$_3372_out0 = v$MUX20_3019_out0[4:0];
assign v$_3372_out1 = v$MUX20_3019_out0[12:8];
assign v$N3_3728_out0 = v$N3_3326_out0;
assign v$N2_680_out0 = v$N2_820_out0;
assign v$N0_1483_out0 = v$_735_out0;
assign v$_1770_out0 = { v$C24_2887_out0,v$_3372_out0 };
assign v$NOTUSE8_4490_out0 = v$_3372_out1;
assign v$N3_4935_out0 = v$N3_3728_out0;
assign v$N1_5023_out0 = v$_500_out0;
assign v$MUX21_779_out0 = v$SEL3_1482_out0 ? v$_1770_out0 : v$MUX20_3019_out0;
assign v$SEL50_2478_out0 = v$N3_4935_out0[20:20];
assign v$N1_2746_out0 = v$N1_5023_out0;
assign v$N2_2836_out0 = v$N2_680_out0;
assign v$N0_3504_out0 = v$N0_1483_out0;
assign v$SEL46_5180_out0 = v$N3_4935_out0[19:10];
assign v$B_83_out0 = v$SEL50_2478_out0;
assign v$SEL6_582_out0 = v$N2_2836_out0[19:19];
assign v$SEL30_1539_out0 = v$N2_2836_out0[20:20];
assign v$N0_1845_out0 = v$N0_3504_out0;
assign v$N1_3180_out0 = v$N1_2746_out0;
assign v$SEL27_3260_out0 = v$N2_2836_out0[18:18];
assign v$SEL29_4444_out0 = v$N2_2836_out0[17:17];
assign v$SEL4_4503_out0 = v$N2_2836_out0[16:7];
assign v$C_4517_out0 = v$SEL46_5180_out0;
assign v$_4766_out0 = v$MUX21_779_out0[8:0];
assign v$_4766_out1 = v$MUX21_779_out0[12:4];
assign v$SEL4_38_out0 = v$C_4517_out0[5:5];
assign v$SEL3_351_out0 = v$N1_3180_out0[16:7];
assign v$SEL25_402_out0 = v$N1_3180_out0[6:6];
assign v$SEL26_466_out0 = v$N1_3180_out0[17:17];
assign v$G4_1353_out0 = ! v$B_83_out0;
assign v$SEL24_1407_out0 = v$C_4517_out0[0:0];
assign v$SEL8_1503_out0 = v$C_4517_out0[4:4];
assign v$SEL30_1613_out0 = v$C_4517_out0[9:9];
assign v$SEL3_1662_out0 = v$C_4517_out0[1:1];
assign v$SEL24_1834_out0 = v$N1_3180_out0[5:5];
assign v$SEL22_2743_out0 = v$N0_1845_out0[6:6];
assign v$SEL1_2795_out0 = v$N0_1845_out0[16:7];
assign v$SEL11_3134_out0 = v$C_4517_out0[3:3];
assign v$SEL28_3406_out0 = v$N1_3180_out0[18:18];
assign v$SEL7_3629_out0 = v$N0_1845_out0[3:0];
assign v$SEL5_3697_out0 = v$N0_1845_out0[4:4];
assign v$SEL2_3922_out0 = v$N1_3180_out0[4:4];
assign v$SEL23_3951_out0 = v$N0_1845_out0[5:5];
assign v$_4008_out0 = { v$C26_1186_out0,v$_4766_out0 };
assign v$SEL21_4308_out0 = v$C_4517_out0[6:6];
assign v$C_4520_out0 = v$SEL4_4503_out0;
assign v$SEL25_4719_out0 = v$C_4517_out0[2:2];
assign v$SEL10_4864_out0 = v$C_4517_out0[8:8];
assign v$A_4989_out0 = v$SEL29_4444_out0;
assign v$A_4998_out0 = v$SEL27_3260_out0;
assign v$SEL14_5214_out0 = v$C_4517_out0[7:7];
assign v$NOTUSE4_5218_out0 = v$_4766_out1;
assign v$C3_27_out0 = v$SEL11_3134_out0;
assign v$SEL4_41_out0 = v$C_4520_out0[5:5];
assign v$B_60_out0 = v$SEL25_402_out0;
assign v$B_79_out0 = v$SEL26_466_out0;
assign v$B_80_out0 = v$SEL2_3922_out0;
assign v$B_87_out0 = v$SEL24_1834_out0;
assign v$B_88_out0 = v$SEL28_3406_out0;
assign v$C2_197_out0 = v$SEL25_4719_out0;
assign v$C9_697_out0 = v$SEL30_1613_out0;
assign v$C0_1107_out0 = v$SEL24_1407_out0;
assign v$C1_1390_out0 = v$SEL3_1662_out0;
assign v$SEL24_1410_out0 = v$C_4520_out0[0:0];
assign v$SEL8_1506_out0 = v$C_4520_out0[4:4];
assign v$SEL30_1616_out0 = v$C_4520_out0[9:9];
assign v$SEL3_1665_out0 = v$C_4520_out0[1:1];
assign v$C8_2448_out0 = v$SEL10_4864_out0;
assign v$MUX18_2657_out0 = v$SEL5_1596_out0 ? v$_4008_out0 : v$MUX21_779_out0;
assign v$G3_2821_out0 = ! v$A_4989_out0;
assign v$G3_2830_out0 = ! v$A_4998_out0;
assign v$SEL11_3137_out0 = v$C_4520_out0[3:3];
assign v$A_3571_out0 = v$SEL3_351_out0;
assign v$B_3843_out0 = v$SEL1_2795_out0;
assign v$C4_4228_out0 = v$SEL8_1503_out0;
assign v$C7_4232_out0 = v$SEL14_5214_out0;
assign v$SEL21_4311_out0 = v$C_4520_out0[6:6];
assign v$C5_4629_out0 = v$SEL4_38_out0;
assign v$SEL25_4722_out0 = v$C_4520_out0[2:2];
assign v$SEL10_4867_out0 = v$C_4520_out0[8:8];
assign v$A_4970_out0 = v$SEL22_2743_out0;
assign v$A_4990_out0 = v$SEL5_3697_out0;
assign v$A_4997_out0 = v$SEL23_3951_out0;
assign v$C6_5170_out0 = v$SEL21_4308_out0;
assign v$SEL14_5217_out0 = v$C_4520_out0[7:7];
assign v$C3_30_out0 = v$SEL11_3137_out0;
assign v$SEL29_99_out0 = v$B_3843_out0[9:9];
assign v$C2_200_out0 = v$SEL25_4722_out0;
assign v$SEL23_587_out0 = v$B_3843_out0[7:7];
assign v$SEL2_606_out0 = v$A_3571_out0[6:6];
assign v$C9_700_out0 = v$SEL30_1616_out0;
assign v$SEL15_833_out0 = v$A_3571_out0[2:2];
assign v$SEL27_920_out0 = v$A_3571_out0[3:3];
assign v$SEL17_995_out0 = v$A_3571_out0[0:0];
assign v$C0_1110_out0 = v$SEL24_1410_out0;
assign v$G4_1330_out0 = ! v$B_60_out0;
assign v$G4_1349_out0 = ! v$B_79_out0;
assign v$G4_1350_out0 = ! v$B_80_out0;
assign v$G4_1357_out0 = ! v$B_87_out0;
assign v$G4_1358_out0 = ! v$B_88_out0;
assign v$C1_1393_out0 = v$SEL3_1665_out0;
assign v$SEL6_1510_out0 = v$B_3843_out0[4:4];
assign v$SEL19_1535_out0 = v$B_3843_out0[2:2];
assign v$SEL26_1766_out0 = v$A_3571_out0[7:7];
assign v$SEL20_1844_out0 = v$B_3843_out0[8:8];
assign v$SEL7_1850_out0 = v$B_3843_out0[0:0];
assign v$SEL16_1898_out0 = v$A_3571_out0[1:1];
assign v$C8_2451_out0 = v$SEL10_4867_out0;
assign v$G1_2536_out0 = v$G3_2821_out0 && v$B_79_out0;
assign v$G1_2545_out0 = v$G3_2830_out0 && v$B_88_out0;
assign v$G3_2802_out0 = ! v$A_4970_out0;
assign v$G3_2822_out0 = ! v$A_4990_out0;
assign v$G3_2829_out0 = ! v$A_4997_out0;
assign v$SEL22_2925_out0 = v$A_3571_out0[8:8];
assign v$SEL13_2984_out0 = v$B_3843_out0[6:6];
assign v$SEL1_3204_out0 = v$A_3571_out0[4:4];
assign v$SEL9_3318_out0 = v$B_3843_out0[1:1];
assign v$_3710_out0 = v$MUX18_2657_out0[10:0];
assign v$_3710_out1 = v$MUX18_2657_out0[12:2];
assign v$SEL12_4142_out0 = v$B_3843_out0[5:5];
assign v$SEL5_4149_out0 = v$A_3571_out0[5:5];
assign v$C4_4231_out0 = v$SEL8_1506_out0;
assign v$C7_4235_out0 = v$SEL14_5217_out0;
assign v$SEL18_4248_out0 = v$B_3843_out0[3:3];
assign v$SEL28_4557_out0 = v$A_3571_out0[9:9];
assign v$C5_4632_out0 = v$SEL4_41_out0;
assign v$C6_5173_out0 = v$SEL21_4311_out0;
assign v$G5_5359_out0 = v$A_4970_out0 && v$B_60_out0;
assign v$G5_5378_out0 = v$A_4989_out0 && v$B_79_out0;
assign v$G5_5379_out0 = v$A_4990_out0 && v$B_80_out0;
assign v$G5_5386_out0 = v$A_4997_out0 && v$B_87_out0;
assign v$G5_5387_out0 = v$A_4998_out0 && v$B_88_out0;
assign v$A6_212_out0 = v$SEL2_606_out0;
assign v$A3_371_out0 = v$SEL27_920_out0;
assign v$C_638_out0 = v$G5_5359_out0;
assign v$C_657_out0 = v$G5_5378_out0;
assign v$C_658_out0 = v$G5_5379_out0;
assign v$C_665_out0 = v$G5_5386_out0;
assign v$C_666_out0 = v$G5_5387_out0;
assign v$B3_879_out0 = v$SEL18_4248_out0;
assign v$A0_916_out0 = v$SEL17_995_out0;
assign v$A9_1283_out0 = v$SEL28_4557_out0;
assign v$B9_1443_out0 = v$SEL29_99_out0;
assign v$A8_1455_out0 = v$SEL22_2925_out0;
assign v$G0_1974_out0 = v$A_4970_out0 && v$G4_1330_out0;
assign v$G0_1993_out0 = v$A_4989_out0 && v$G4_1349_out0;
assign v$G0_1994_out0 = v$A_4990_out0 && v$G4_1350_out0;
assign v$G0_2001_out0 = v$A_4997_out0 && v$G4_1357_out0;
assign v$G0_2002_out0 = v$A_4998_out0 && v$G4_1358_out0;
assign v$A4_2223_out0 = v$SEL1_3204_out0;
assign v$B4_2252_out0 = v$SEL6_1510_out0;
assign v$G1_2517_out0 = v$G3_2802_out0 && v$B_60_out0;
assign v$G1_2537_out0 = v$G3_2822_out0 && v$B_80_out0;
assign v$G1_2544_out0 = v$G3_2829_out0 && v$B_87_out0;
assign v$B2_2648_out0 = v$SEL19_1535_out0;
assign v$B6_2665_out0 = v$SEL13_2984_out0;
assign v$A2_2731_out0 = v$SEL15_833_out0;
assign v$_2837_out0 = { v$C22_3079_out0,v$_3710_out0 };
assign v$B8_3057_out0 = v$SEL20_1844_out0;
assign v$B1_3238_out0 = v$SEL9_3318_out0;
assign v$A1_3823_out0 = v$SEL16_1898_out0;
assign v$B7_3921_out0 = v$SEL23_587_out0;
assign v$B5_4007_out0 = v$SEL12_4142_out0;
assign v$A7_4166_out0 = v$SEL26_1766_out0;
assign v$B0_4343_out0 = v$SEL7_1850_out0;
assign v$NOTUSE2_4541_out0 = v$_3710_out1;
assign v$A5_4741_out0 = v$SEL5_4149_out0;
assign {v$A4_345_out1,v$A4_345_out0 } = v$B1_3238_out0 + v$C1_1393_out0 + v$A1_3823_out0;
assign v$G2_429_out0 = v$G0_1974_out0 || v$G1_2517_out0;
assign v$G2_448_out0 = v$G0_1993_out0 || v$G1_2536_out0;
assign v$G2_449_out0 = v$G0_1994_out0 || v$G1_2537_out0;
assign v$G2_456_out0 = v$G0_2001_out0 || v$G1_2544_out0;
assign v$G2_457_out0 = v$G0_2002_out0 || v$G1_2545_out0;
assign {v$A1_1302_out1,v$A1_1302_out0 } = v$B4_2252_out0 + v$C4_4231_out0 + v$A4_2223_out0;
assign v$MUX19_1397_out0 = v$SEL2_4934_out0 ? v$_2837_out0 : v$MUX18_2657_out0;
assign {v$A8_1631_out1,v$A8_1631_out0 } = v$B8_3057_out0 + v$C8_2451_out0 + v$A8_1455_out0;
assign {v$A6_1659_out1,v$A6_1659_out0 } = v$B6_2665_out0 + v$C6_5173_out0 + v$A6_212_out0;
assign v$_1779_out0 = { v$C_665_out0,v$C_638_out0 };
assign v$_2129_out0 = { v$C_657_out0,v$C_666_out0 };
assign {v$A10_3268_out1,v$A10_3268_out0 } = v$B9_1443_out0 + v$C9_700_out0 + v$A9_1283_out0;
assign v$_3583_out0 = { v$C1_2666_out0,v$C_658_out0 };
assign {v$A7_3671_out1,v$A7_3671_out0 } = v$B0_4343_out0 + v$C0_1110_out0 + v$A0_916_out0;
assign {v$A9_3766_out1,v$A9_3766_out0 } = v$B5_4007_out0 + v$C5_4632_out0 + v$A5_4741_out0;
assign {v$A2_4331_out1,v$A2_4331_out0 } = v$B3_879_out0 + v$C3_30_out0 + v$A3_371_out0;
assign {v$A5_4642_out1,v$A5_4642_out0 } = v$B2_2648_out0 + v$C2_200_out0 + v$A2_2731_out0;
assign {v$A3_5329_out1,v$A3_5329_out0 } = v$B7_3921_out0 + v$C7_4235_out0 + v$A7_4166_out0;
assign v$S12_103_out0 = v$A5_4642_out1;
assign v$S19_571_out0 = v$A10_3268_out1;
assign v$S14_670_out0 = v$A1_1302_out1;
assign v$S13_854_out0 = v$A2_4331_out1;
assign v$S07_889_out0 = v$A3_5329_out0;
assign v$S10_941_out0 = v$A7_3671_out1;
assign v$S01_1064_out0 = v$A4_345_out0;
assign v$S08_1592_out0 = v$A8_1631_out0;
assign v$_1811_out0 = v$MUX19_1397_out0[11:0];
assign v$_1811_out1 = v$MUX19_1397_out0[12:1];
assign v$S09_1939_out0 = v$A10_3268_out0;
assign v$_2068_out0 = { v$_3583_out0,v$_1779_out0 };
assign v$S04_2281_out0 = v$A1_1302_out0;
assign v$S18_2439_out0 = v$A8_1631_out1;
assign v$S03_2847_out0 = v$A2_4331_out0;
assign v$S06_3114_out0 = v$A6_1659_out0;
assign v$S11_3143_out0 = v$A4_345_out1;
assign v$S15_3219_out0 = v$A9_3766_out1;
assign v$S02_3393_out0 = v$A5_4642_out0;
assign v$S17_4093_out0 = v$A3_5329_out1;
assign v$S_4175_out0 = v$G2_429_out0;
assign v$S_4194_out0 = v$G2_448_out0;
assign v$S_4195_out0 = v$G2_449_out0;
assign v$S_4202_out0 = v$G2_456_out0;
assign v$S_4203_out0 = v$G2_457_out0;
assign v$S00_4442_out0 = v$A7_3671_out0;
assign v$S16_4697_out0 = v$A6_1659_out1;
assign v$S05_4889_out0 = v$A9_3766_out0;
assign v$_177_out0 = { v$S08_1592_out0,v$S09_1939_out0 };
assign v$_239_out0 = { v$S18_2439_out0,v$S19_571_out0 };
assign v$_946_out0 = { v$S02_3393_out0,v$S03_2847_out0 };
assign v$_1166_out0 = { v$S00_4442_out0,v$S01_1064_out0 };
assign v$_1797_out0 = { v$S_4203_out0,v$SEL6_582_out0 };
assign v$_1891_out0 = { v$S16_4697_out0,v$S17_4093_out0 };
assign v$_2737_out0 = { v$S10_941_out0,v$S11_3143_out0 };
assign v$_2939_out0 = { v$C23_979_out0,v$_1811_out0 };
assign v$_3035_out0 = { v$SEL7_3629_out0,v$S_4195_out0 };
assign v$_3110_out0 = { v$S14_670_out0,v$S15_3219_out0 };
assign v$_3363_out0 = { v$S_4202_out0,v$S_4175_out0 };
assign v$_3578_out0 = { v$S06_3114_out0,v$S07_889_out0 };
assign v$_3817_out0 = { v$S12_103_out0,v$S13_854_out0 };
assign v$NOTUSE1_4377_out0 = v$_1811_out1;
assign v$_4881_out0 = { v$S04_2281_out0,v$S05_4889_out0 };
assign v$_1423_out0 = { v$_2737_out0,v$_3817_out0 };
assign v$_1673_out0 = { v$_4881_out0,v$_3578_out0 };
assign v$MUX17_1753_out0 = v$SEL1_4771_out0 ? v$_2939_out0 : v$MUX19_1397_out0;
assign v$_2020_out0 = { v$_3110_out0,v$_1891_out0 };
assign v$_2076_out0 = { v$_1166_out0,v$_946_out0 };
assign v$_690_out0 = { v$_1673_out0,v$_177_out0 };
assign v$OUTPUT_3581_out0 = v$MUX17_1753_out0;
assign v$_4059_out0 = { v$_2020_out0,v$_239_out0 };
assign v$_3041_out0 = { v$_1423_out0,v$_4059_out0 };
assign v$_3611_out0 = { v$_2076_out0,v$_690_out0 };
assign v$_5259_out0 = v$OUTPUT_3581_out0[1:0];
assign v$_5259_out1 = v$OUTPUT_3581_out0[12:11];
assign v$_1927_out0 = v$_5259_out1[9:0];
assign v$_1927_out1 = v$_5259_out1[10:1];
assign v$ROUNDING_3068_out0 = v$_5259_out0;
assign v$S1_4208_out0 = v$_3611_out0;
assign v$S2_4318_out0 = v$_3041_out0;
assign v$NEWFRAC_608_out0 = v$_1927_out0;
assign v$_3536_out0 = { v$S2_4318_out0,v$_2129_out0 };
assign v$INT_3598_out0 = v$_1927_out1;
assign v$_4536_out0 = { v$S1_4208_out0,v$S_4194_out0 };
assign v$_2755_out0 = { v$_3536_out0,v$SEL30_1539_out0 };
assign v$_3560_out0 = { v$_3363_out0,v$_4536_out0 };
assign v$_3784_out0 = { v$NEWFRAC_608_out0,v$NEWEXPO_4492_out0 };
assign v$_980_out0 = { v$_2068_out0,v$_2755_out0 };
assign v$_2774_out0 = { v$_3560_out0,v$_1797_out0 };
assign v$fpmerge_5196_out0 = { v$_3784_out0,v$NEWSIGN_3096_out0 };
assign v$_3589_out0 = { v$_3035_out0,v$_2774_out0 };
assign v$1_4825_out0 = v$_980_out0;
assign v$SEL32_36_out0 = v$1_4825_out0[7:7];
assign v$SEL33_1035_out0 = v$1_4825_out0[8:8];
assign v$SEL43_1956_out0 = v$1_4825_out0[5:5];
assign v$SEL49_2881_out0 = v$1_4825_out0[20:20];
assign v$SEL36_3144_out0 = v$1_4825_out0[6:6];
assign v$SEL40_4711_out0 = v$1_4825_out0[9:9];
assign v$0_5061_out0 = v$_3589_out0;
assign v$SEL31_5225_out0 = v$1_4825_out0[19:10];
assign v$B_78_out0 = v$SEL40_4711_out0;
assign v$B_81_out0 = v$SEL33_1035_out0;
assign v$B_82_out0 = v$SEL36_3144_out0;
assign v$B_84_out0 = v$SEL32_36_out0;
assign v$B_86_out0 = v$SEL43_1956_out0;
assign v$SEL38_465_out0 = v$0_5061_out0[19:10];
assign v$SEL41_975_out0 = v$0_5061_out0[4:0];
assign v$SEL47_1719_out0 = v$0_5061_out0[8:8];
assign v$SEL42_2134_out0 = v$0_5061_out0[5:5];
assign v$SEL44_2612_out0 = v$0_5061_out0[6:6];
assign v$SEL37_2633_out0 = v$0_5061_out0[7:7];
assign v$A_3568_out0 = v$SEL31_5225_out0;
assign v$SEL48_3948_out0 = v$0_5061_out0[9:9];
assign v$A_4993_out0 = v$SEL49_2881_out0;
assign v$SEL2_603_out0 = v$A_3568_out0[6:6];
assign v$SEL15_830_out0 = v$A_3568_out0[2:2];
assign v$SEL27_917_out0 = v$A_3568_out0[3:3];
assign v$SEL17_992_out0 = v$A_3568_out0[0:0];
assign v$G4_1348_out0 = ! v$B_78_out0;
assign v$G4_1351_out0 = ! v$B_81_out0;
assign v$G4_1352_out0 = ! v$B_82_out0;
assign v$G4_1354_out0 = ! v$B_84_out0;
assign v$G4_1356_out0 = ! v$B_86_out0;
assign v$SEL26_1763_out0 = v$A_3568_out0[7:7];
assign v$SEL16_1895_out0 = v$A_3568_out0[1:1];
assign v$G0_1997_out0 = v$A_4993_out0 && v$G4_1353_out0;
assign v$G3_2825_out0 = ! v$A_4993_out0;
assign v$SEL22_2922_out0 = v$A_3568_out0[8:8];
assign v$SEL1_3201_out0 = v$A_3568_out0[4:4];
assign v$B_3840_out0 = v$SEL38_465_out0;
assign v$SEL5_4146_out0 = v$A_3568_out0[5:5];
assign v$SEL28_4554_out0 = v$A_3568_out0[9:9];
assign v$A_4988_out0 = v$SEL48_3948_out0;
assign v$A_4991_out0 = v$SEL47_1719_out0;
assign v$A_4992_out0 = v$SEL44_2612_out0;
assign v$A_4994_out0 = v$SEL37_2633_out0;
assign v$A_4996_out0 = v$SEL42_2134_out0;
assign v$G5_5382_out0 = v$A_4993_out0 && v$B_83_out0;
assign v$SEL29_96_out0 = v$B_3840_out0[9:9];
assign v$A6_209_out0 = v$SEL2_603_out0;
assign v$A3_368_out0 = v$SEL27_917_out0;
assign v$SEL23_584_out0 = v$B_3840_out0[7:7];
assign v$C_661_out0 = v$G5_5382_out0;
assign v$A0_913_out0 = v$SEL17_992_out0;
assign v$A9_1280_out0 = v$SEL28_4554_out0;
assign v$A8_1452_out0 = v$SEL22_2922_out0;
assign v$SEL6_1507_out0 = v$B_3840_out0[4:4];
assign v$SEL19_1532_out0 = v$B_3840_out0[2:2];
assign v$SEL20_1841_out0 = v$B_3840_out0[8:8];
assign v$SEL7_1847_out0 = v$B_3840_out0[0:0];
assign v$G0_1992_out0 = v$A_4988_out0 && v$G4_1348_out0;
assign v$G0_1995_out0 = v$A_4991_out0 && v$G4_1351_out0;
assign v$G0_1996_out0 = v$A_4992_out0 && v$G4_1352_out0;
assign v$G0_1998_out0 = v$A_4994_out0 && v$G4_1354_out0;
assign v$G0_2000_out0 = v$A_4996_out0 && v$G4_1356_out0;
assign v$A4_2220_out0 = v$SEL1_3201_out0;
assign v$G1_2540_out0 = v$G3_2825_out0 && v$B_83_out0;
assign v$A2_2728_out0 = v$SEL15_830_out0;
assign v$G3_2820_out0 = ! v$A_4988_out0;
assign v$G3_2823_out0 = ! v$A_4991_out0;
assign v$G3_2824_out0 = ! v$A_4992_out0;
assign v$G3_2826_out0 = ! v$A_4994_out0;
assign v$G3_2828_out0 = ! v$A_4996_out0;
assign v$SEL13_2981_out0 = v$B_3840_out0[6:6];
assign v$SEL9_3315_out0 = v$B_3840_out0[1:1];
assign v$A1_3820_out0 = v$SEL16_1895_out0;
assign v$SEL12_4139_out0 = v$B_3840_out0[5:5];
assign v$A7_4163_out0 = v$SEL26_1763_out0;
assign v$SEL18_4245_out0 = v$B_3840_out0[3:3];
assign v$A5_4738_out0 = v$SEL5_4146_out0;
assign v$G5_5377_out0 = v$A_4988_out0 && v$B_78_out0;
assign v$G5_5380_out0 = v$A_4991_out0 && v$B_81_out0;
assign v$G5_5381_out0 = v$A_4992_out0 && v$B_82_out0;
assign v$G5_5383_out0 = v$A_4994_out0 && v$B_84_out0;
assign v$G5_5385_out0 = v$A_4996_out0 && v$B_86_out0;
assign v$G2_452_out0 = v$G0_1997_out0 || v$G1_2540_out0;
assign v$C_656_out0 = v$G5_5377_out0;
assign v$C_659_out0 = v$G5_5380_out0;
assign v$C_660_out0 = v$G5_5381_out0;
assign v$C_662_out0 = v$G5_5383_out0;
assign v$C_664_out0 = v$G5_5385_out0;
assign v$B3_876_out0 = v$SEL18_4245_out0;
assign v$B9_1440_out0 = v$SEL29_96_out0;
assign v$B4_2249_out0 = v$SEL6_1507_out0;
assign v$G1_2535_out0 = v$G3_2820_out0 && v$B_78_out0;
assign v$G1_2538_out0 = v$G3_2823_out0 && v$B_81_out0;
assign v$G1_2539_out0 = v$G3_2824_out0 && v$B_82_out0;
assign v$G1_2541_out0 = v$G3_2826_out0 && v$B_84_out0;
assign v$G1_2543_out0 = v$G3_2828_out0 && v$B_86_out0;
assign v$B2_2645_out0 = v$SEL19_1532_out0;
assign v$B6_2662_out0 = v$SEL13_2981_out0;
assign v$B8_3054_out0 = v$SEL20_1841_out0;
assign v$B1_3235_out0 = v$SEL9_3315_out0;
assign v$B7_3918_out0 = v$SEL23_584_out0;
assign v$B5_4004_out0 = v$SEL12_4139_out0;
assign v$B0_4340_out0 = v$SEL7_1847_out0;
assign {v$A4_342_out1,v$A4_342_out0 } = v$B1_3235_out0 + v$C1_1390_out0 + v$A1_3820_out0;
assign v$G2_447_out0 = v$G0_1992_out0 || v$G1_2535_out0;
assign v$G2_450_out0 = v$G0_1995_out0 || v$G1_2538_out0;
assign v$G2_451_out0 = v$G0_1996_out0 || v$G1_2539_out0;
assign v$G2_453_out0 = v$G0_1998_out0 || v$G1_2541_out0;
assign v$G2_455_out0 = v$G0_2000_out0 || v$G1_2543_out0;
assign {v$A1_1299_out1,v$A1_1299_out0 } = v$B4_2249_out0 + v$C4_4228_out0 + v$A4_2220_out0;
assign {v$A8_1628_out1,v$A8_1628_out0 } = v$B8_3054_out0 + v$C8_2448_out0 + v$A8_1452_out0;
assign {v$A6_1656_out1,v$A6_1656_out0 } = v$B6_2662_out0 + v$C6_5170_out0 + v$A6_209_out0;
assign v$_1903_out0 = { v$C5_4278_out0,v$C_664_out0 };
assign v$_2694_out0 = { v$C_660_out0,v$C_662_out0 };
assign {v$A10_3265_out1,v$A10_3265_out0 } = v$B9_1440_out0 + v$C9_697_out0 + v$A9_1280_out0;
assign {v$A7_3668_out1,v$A7_3668_out0 } = v$B0_4340_out0 + v$C0_1107_out0 + v$A0_913_out0;
assign {v$A9_3763_out1,v$A9_3763_out0 } = v$B5_4004_out0 + v$C5_4629_out0 + v$A5_4738_out0;
assign v$_4073_out0 = { v$C_659_out0,v$C_656_out0 };
assign v$S_4198_out0 = v$G2_452_out0;
assign {v$A2_4328_out1,v$A2_4328_out0 } = v$B3_876_out0 + v$C3_27_out0 + v$A3_368_out0;
assign {v$A5_4639_out1,v$A5_4639_out0 } = v$B2_2645_out0 + v$C2_197_out0 + v$A2_2728_out0;
assign {v$A3_5326_out1,v$A3_5326_out0 } = v$B7_3918_out0 + v$C7_4232_out0 + v$A7_4163_out0;
assign v$S12_100_out0 = v$A5_4639_out1;
assign v$S19_568_out0 = v$A10_3265_out1;
assign v$S14_667_out0 = v$A1_1299_out1;
assign v$S13_851_out0 = v$A2_4328_out1;
assign v$S07_886_out0 = v$A3_5326_out0;
assign v$S10_938_out0 = v$A7_3668_out1;
assign v$S01_1061_out0 = v$A4_342_out0;
assign v$S08_1589_out0 = v$A8_1628_out0;
assign v$S09_1936_out0 = v$A10_3265_out0;
assign v$S04_2278_out0 = v$A1_1299_out0;
assign v$S18_2436_out0 = v$A8_1628_out1;
assign v$S03_2844_out0 = v$A2_4328_out0;
assign v$S06_3111_out0 = v$A6_1656_out0;
assign v$S11_3140_out0 = v$A4_342_out1;
assign v$S15_3216_out0 = v$A9_3763_out1;
assign v$S02_3390_out0 = v$A5_4639_out0;
assign v$_4016_out0 = { v$_1903_out0,v$_2694_out0 };
assign v$S17_4090_out0 = v$A3_5326_out1;
assign v$S_4193_out0 = v$G2_447_out0;
assign v$S_4196_out0 = v$G2_450_out0;
assign v$S_4197_out0 = v$G2_451_out0;
assign v$S_4199_out0 = v$G2_453_out0;
assign v$S_4201_out0 = v$G2_455_out0;
assign v$S00_4439_out0 = v$A7_3668_out0;
assign v$S16_4694_out0 = v$A6_1656_out1;
assign v$S05_4886_out0 = v$A9_3763_out0;
assign v$_174_out0 = { v$S08_1589_out0,v$S09_1936_out0 };
assign v$_236_out0 = { v$S18_2436_out0,v$S19_568_out0 };
assign v$_498_out0 = { v$S_4196_out0,v$S_4193_out0 };
assign v$_943_out0 = { v$S02_3390_out0,v$S03_2844_out0 };
assign v$_1163_out0 = { v$S00_4439_out0,v$S01_1061_out0 };
assign v$_1888_out0 = { v$S16_4694_out0,v$S17_4090_out0 };
assign v$_1965_out0 = { v$S_4197_out0,v$S_4199_out0 };
assign v$_2734_out0 = { v$S10_938_out0,v$S11_3140_out0 };
assign v$_3107_out0 = { v$S14_667_out0,v$S15_3216_out0 };
assign v$_3575_out0 = { v$S06_3111_out0,v$S07_886_out0 };
assign v$_3814_out0 = { v$S12_100_out0,v$S13_851_out0 };
assign v$_4749_out0 = { v$SEL41_975_out0,v$S_4201_out0 };
assign v$_4878_out0 = { v$S04_2278_out0,v$S05_4886_out0 };
assign v$_316_out0 = { v$_1965_out0,v$_498_out0 };
assign v$_1420_out0 = { v$_2734_out0,v$_3814_out0 };
assign v$_1670_out0 = { v$_4878_out0,v$_3575_out0 };
assign v$_2017_out0 = { v$_3107_out0,v$_1888_out0 };
assign v$_2073_out0 = { v$_1163_out0,v$_943_out0 };
assign v$_687_out0 = { v$_1670_out0,v$_174_out0 };
assign v$_4056_out0 = { v$_2017_out0,v$_236_out0 };
assign v$_3038_out0 = { v$_1420_out0,v$_4056_out0 };
assign v$_3608_out0 = { v$_2073_out0,v$_687_out0 };
assign v$S1_4205_out0 = v$_3608_out0;
assign v$S2_4315_out0 = v$_3038_out0;
assign v$_1786_out0 = { v$S2_4315_out0,v$C_661_out0 };
assign v$_3580_out0 = { v$S1_4205_out0,v$S_4198_out0 };
assign v$_1900_out0 = { v$_316_out0,v$_3580_out0 };
assign v$_4730_out0 = { v$_4073_out0,v$_1786_out0 };
assign v$_1264_out0 = { v$_4749_out0,v$_1900_out0 };
assign v$_1417_out0 = { v$_4016_out0,v$_4730_out0 };
assign v$00_1369_out0 = v$_1264_out0;
assign v$11_2653_out0 = v$_1417_out0;
assign v$SEL52_1439_out0 = v$11_2653_out0[20:6];
assign v$SEL53_3630_out0 = v$00_1369_out0[20:6];
assign v$SEL54_4089_out0 = v$11_2653_out0[21:21];
assign v$SEL51_4277_out0 = v$00_1369_out0[5:0];
assign v$B_85_out0 = v$SEL54_4089_out0;
assign {v$A1_794_out1,v$A1_794_out0 } = v$SEL52_1439_out0 + v$SEL53_3630_out0 + v$C6_702_out0;
assign v$G4_1355_out0 = ! v$B_85_out0;
assign v$_4209_out0 = { v$SEL51_4277_out0,v$A1_794_out0 };
assign v$A_4995_out0 = v$A1_794_out1;
assign v$G0_1999_out0 = v$A_4995_out0 && v$G4_1355_out0;
assign v$G3_2827_out0 = ! v$A_4995_out0;
assign v$G5_5384_out0 = v$A_4995_out0 && v$B_85_out0;
assign v$C_663_out0 = v$G5_5384_out0;
assign v$G1_2542_out0 = v$G3_2827_out0 && v$B_85_out0;
assign v$G2_454_out0 = v$G0_1999_out0 || v$G1_2542_out0;
assign v$X_1263_out0 = v$C_663_out0;
assign v$S_4200_out0 = v$G2_454_out0;
assign v$_2181_out0 = { v$_4209_out0,v$S_4200_out0 };
assign v$OUTPUT_1902_out0 = v$_2181_out0;
assign v$FRAC_1303_out0 = v$OUTPUT_1902_out0;
assign v$IN_1444_out0 = v$OUTPUT_1902_out0;
assign v$INPUT_2972_out0 = v$OUTPUT_1902_out0;
assign v$FRAC22_4051_out0 = v$OUTPUT_1902_out0;
assign v$SEL2_817_out0 = v$FRAC_1303_out0[21:20];
assign v$_2006_out0 = v$INPUT_2972_out0[20:0];
assign v$_2006_out1 = v$INPUT_2972_out0[21:1];
assign v$SEL1_2548_out0 = v$FRAC_1303_out0[21:21];
assign v$_2865_out0 = v$IN_1444_out0[20:0];
assign v$_2865_out1 = v$IN_1444_out0[21:1];
assign v$_3335_out0 = v$FRAC_1303_out0[0:0];
assign v$_3335_out1 = v$FRAC_1303_out0[21:21];
assign v$IN1_3927_out0 = v$FRAC22_4051_out0;
assign v$X1_1220_out0 = v$_3335_out0;
assign v$_2516_out0 = v$_2006_out0[7:0];
assign v$_2516_out1 = v$_2006_out0[20:13];
assign v$_2849_out0 = { v$_3335_out1,v$C2_4034_out0 };
assign v$_2987_out0 = v$_2865_out0[19:0];
assign v$_2987_out1 = v$_2865_out0[20:1];
assign v$SEL2_3384_out0 = v$IN1_3927_out0[21:21];
assign v$EQ2_3619_out0 = v$SEL2_817_out0 == 2'h1;
assign v$NOTUSEMSB_4611_out0 = v$_2865_out1;
assign v$RIGHTSHIFT_4693_out0 = v$SEL1_2548_out0;
assign v$MSB_4908_out0 = v$_2006_out1;
assign v$_5096_out0 = v$IN1_3927_out0[0:0];
assign v$_5096_out1 = v$IN1_3927_out0[21:21];
assign v$EXPONOCHANGE_278_out0 = v$EQ2_3619_out0;
assign v$_416_out0 = { v$C2_23_out0,v$_2987_out0 };
assign v$X_530_out0 = v$_2987_out1;
assign v$MSB_1458_out0 = v$SEL2_3384_out0;
assign v$_2375_out0 = { v$_5096_out1,v$C1_2702_out0 };
assign {v$A1_2427_out1,v$A1_2427_out0 } = v$SEL4_676_out0 + v$C1_3138_out0 + v$RIGHTSHIFT_4693_out0;
assign v$INPUT_3071_out0 = v$_2516_out1;
assign v$INPUT_3072_out0 = v$_2516_out0;
assign v$X5_4793_out0 = v$_5096_out0;
assign v$MUX2_5410_out0 = v$RIGHTSHIFT_4693_out0 ? v$_2849_out0 : v$FRAC_1303_out0;
assign v$SEL18_24_out0 = v$INPUT_3071_out0[3:3];
assign v$SEL18_25_out0 = v$INPUT_3072_out0[3:3];
assign v$NEWFRAC_249_out0 = v$MUX2_5410_out0;
assign v$SEL5_266_out0 = v$INPUT_3071_out0[10:10];
assign v$SEL15_467_out0 = v$INPUT_3071_out0[4:4];
assign v$SEL15_468_out0 = v$INPUT_3072_out0[4:4];
assign v$X_759_out0 = v$A1_2427_out1;
assign v$MUX2_974_out0 = v$1_4568_out0 ? v$_2375_out0 : v$IN1_3927_out0;
assign v$SEL14_1153_out0 = v$INPUT_3071_out0[7:7];
assign v$SEL14_1154_out0 = v$INPUT_3072_out0[7:7];
assign v$SEL12_1173_out0 = v$INPUT_3071_out0[12:12];
assign v$SEL7_1405_out0 = v$INPUT_3071_out0[8:8];
assign v$SEL6_1560_out0 = v$INPUT_3071_out0[9:9];
assign v$SEL21_2091_out0 = v$INPUT_3071_out0[0:0];
assign v$SEL21_2092_out0 = v$INPUT_3072_out0[0:0];
assign v$MUX1_2143_out0 = v$EXPONOCHANGE_278_out0 ? v$SEL4_676_out0 : v$A1_2427_out0;
assign v$SEL20_2270_out0 = v$INPUT_3071_out0[1:1];
assign v$SEL20_2271_out0 = v$INPUT_3072_out0[1:1];
assign v$SEL13_3455_out0 = v$INPUT_3071_out0[6:6];
assign v$SEL13_3456_out0 = v$INPUT_3072_out0[6:6];
assign v$SEL17_3944_out0 = v$INPUT_3071_out0[2:2];
assign v$SEL17_3945_out0 = v$INPUT_3072_out0[2:2];
assign v$SEL16_4038_out0 = v$INPUT_3071_out0[5:5];
assign v$SEL16_4039_out0 = v$INPUT_3072_out0[5:5];
assign v$SEL1_4767_out0 = v$INPUT_3071_out0[11:11];
assign v$G52_301_out0 = ! v$SEL15_467_out0;
assign v$G52_302_out0 = ! v$SEL15_468_out0;
assign v$G66_557_out0 = ! v$SEL21_2091_out0;
assign v$G46_559_out0 = ! v$SEL13_3455_out0;
assign v$G46_560_out0 = ! v$SEL13_3456_out0;
assign v$SEL5_701_out0 = v$MUX1_2143_out0[5:5];
assign v$G19_786_out0 = ! v$SEL5_266_out0;
assign v$G17_1082_out0 = ! v$SEL1_4767_out0;
assign v$G39_1318_out0 = ! v$SEL12_1173_out0;
assign v$NEWFRAC1011_2046_out0 = v$NEWFRAC_249_out0;
assign v$_2097_out0 = v$MUX2_974_out0[1:0];
assign v$_2097_out1 = v$MUX2_974_out0[21:20];
assign v$G40_2289_out0 = ! v$SEL7_1405_out0;
assign v$G45_2791_out0 = ! v$SEL14_1153_out0;
assign v$G45_2792_out0 = ! v$SEL14_1154_out0;
assign v$SEL6_3327_out0 = v$MUX1_2143_out0[4:0];
assign v$G22_3336_out0 = ! v$SEL6_1560_out0;
assign v$G51_3595_out0 = ! v$SEL16_4038_out0;
assign v$G51_3596_out0 = ! v$SEL16_4039_out0;
assign v$G58_4583_out0 = ! v$SEL17_3944_out0;
assign v$G58_4584_out0 = ! v$SEL17_3945_out0;
assign v$G57_4883_out0 = ! v$SEL18_24_out0;
assign v$G57_4884_out0 = ! v$SEL18_25_out0;
assign v$G62_4941_out0 = ! v$SEL20_2270_out0;
assign v$G62_4942_out0 = ! v$SEL20_2271_out0;
assign v$12_5202_out0 = v$SEL12_1173_out0;
assign v$MUX13_849_out0 = v$12_5202_out0 ? v$C2_4459_out0 : v$C1_2298_out0;
assign v$G18_2013_out0 = v$G17_1082_out0 && v$G39_1318_out0;
assign v$X8_2515_out0 = v$_2097_out0;
assign v$OVERFLOW_2597_out0 = v$SEL5_701_out0;
assign v$G6_3367_out0 = v$SEL1_4767_out0 && v$G39_1318_out0;
assign v$NEWEXPO_4385_out0 = v$SEL6_3327_out0;
assign v$_4616_out0 = { v$_2097_out1,v$C8_338_out0 };
assign v$G20_318_out0 = v$SEL5_266_out0 && v$G18_2013_out0;
assign v$MUX8_349_out0 = v$2_3042_out0 ? v$_4616_out0 : v$MUX2_974_out0;
assign v$G23_1484_out0 = v$G19_786_out0 && v$G18_2013_out0;
assign v$OVERFLOW1_4085_out0 = v$OVERFLOW_2597_out0;
assign v$11_4305_out0 = v$G6_3367_out0;
assign v$NEWEXPO1011_4381_out0 = v$NEWEXPO_4385_out0;
assign v$10_548_out0 = v$G20_318_out0;
assign v$G26_818_out0 = v$G22_3336_out0 && v$G23_1484_out0;
assign v$_972_out0 = v$MUX8_349_out0[2:0];
assign v$_972_out1 = v$MUX8_349_out0[21:19];
assign v$G21_1800_out0 = v$SEL6_1560_out0 && v$G23_1484_out0;
assign v$MUX9_3445_out0 = v$11_4305_out0 ? v$C3_5357_out0 : v$MUX13_849_out0;
assign v$_5136_out0 = { v$12_5202_out0,v$11_4305_out0 };
assign v$X6_673_out0 = v$_972_out0;
assign v$_1735_out0 = { v$_972_out1,v$C4_2077_out0 };
assign v$9_2615_out0 = v$G21_1800_out0;
assign v$G24_2700_out0 = v$SEL7_1405_out0 && v$G26_818_out0;
assign v$G42_2707_out0 = v$G40_2289_out0 && v$G26_818_out0;
assign v$MUX12_3905_out0 = v$10_548_out0 ? v$C4_1031_out0 : v$MUX9_3445_out0;
assign v$MUX10_589_out0 = v$9_2615_out0 ? v$C5_4464_out0 : v$MUX12_3905_out0;
assign v$_1069_out0 = { v$10_548_out0,v$9_2615_out0 };
assign v$G41_1466_out0 = v$G45_2791_out0 && v$G42_2707_out0;
assign v$8_1972_out0 = v$G24_2700_out0;
assign v$G43_2433_out0 = v$SEL14_1153_out0 && v$G42_2707_out0;
assign v$MUX11_3385_out0 = v$3_490_out0 ? v$_1735_out0 : v$MUX8_349_out0;
assign v$_365_out0 = v$MUX11_3385_out0[3:0];
assign v$_365_out1 = v$MUX11_3385_out0[21:18];
assign v$MUX11_1881_out0 = v$8_1972_out0 ? v$C6_4823_out0 : v$MUX10_589_out0;
assign v$G48_2725_out0 = v$G46_559_out0 && v$G41_1466_out0;
assign v$G44_3209_out0 = v$SEL13_3455_out0 && v$G41_1466_out0;
assign v$_3599_out0 = { v$_5136_out0,v$_1069_out0 };
assign v$7_4951_out0 = v$G43_2433_out0;
assign v$_58_out0 = { v$_365_out1,v$C10_1253_out0 };
assign v$_1746_out0 = { v$8_1972_out0,v$7_4951_out0 };
assign v$MUX8_2408_out0 = v$7_4951_out0 ? v$C7_1908_out0 : v$MUX11_1881_out0;
assign v$X11_3193_out0 = v$_365_out0;
assign v$G49_3412_out0 = v$SEL16_4038_out0 && v$G48_2725_out0;
assign v$6_3495_out0 = v$G44_3209_out0;
assign v$G47_4373_out0 = v$G51_3595_out0 && v$G48_2725_out0;
assign v$G50_246_out0 = v$SEL15_467_out0 && v$G47_4373_out0;
assign v$G54_2008_out0 = v$G52_301_out0 && v$G47_4373_out0;
assign v$MUX6_3118_out0 = v$6_3495_out0 ? v$C8_2634_out0 : v$MUX8_2408_out0;
assign v$MUX9_3900_out0 = v$4_718_out0 ? v$_58_out0 : v$MUX11_3385_out0;
assign v$5_4219_out0 = v$G49_3412_out0;
assign v$_1046_out0 = v$MUX9_3900_out0[4:0];
assign v$_1046_out1 = v$MUX9_3900_out0[21:17];
assign v$4_1200_out0 = v$G50_246_out0;
assign v$MUX5_1751_out0 = v$5_4219_out0 ? v$C9_2796_out0 : v$MUX6_3118_out0;
assign v$G53_2295_out0 = v$G57_4883_out0 && v$G54_2008_out0;
assign v$G55_3407_out0 = v$SEL18_24_out0 && v$G54_2008_out0;
assign v$_4788_out0 = { v$6_3495_out0,v$5_4219_out0 };
assign v$MUX7_525_out0 = v$4_1200_out0 ? v$C10_1968_out0 : v$MUX5_1751_out0;
assign v$_716_out0 = { v$_1046_out1,v$C6_2426_out0 };
assign v$G56_2854_out0 = v$SEL17_3944_out0 && v$G53_2295_out0;
assign v$_3120_out0 = { v$_1746_out0,v$_4788_out0 };
assign v$X2_3685_out0 = v$_1046_out0;
assign v$3_4626_out0 = v$G55_3407_out0;
assign v$G60_5426_out0 = v$G58_4583_out0 && v$G53_2295_out0;
assign v$_20_out0 = { v$4_1200_out0,v$3_4626_out0 };
assign v$MUX4_725_out0 = v$3_4626_out0 ? v$C11_3342_out0 : v$MUX7_525_out0;
assign v$G63_821_out0 = v$G62_4941_out0 && v$G60_5426_out0;
assign v$_2315_out0 = { v$_3599_out0,v$_3120_out0 };
assign v$2_2917_out0 = v$G56_2854_out0;
assign v$G61_3941_out0 = v$SEL20_2270_out0 && v$G60_5426_out0;
assign v$MUX7_4758_out0 = v$5_2475_out0 ? v$_716_out0 : v$MUX9_3900_out0;
assign v$G65_130_out0 = v$G66_557_out0 && v$G63_821_out0;
assign v$G64_2688_out0 = v$G63_821_out0 && v$SEL21_2091_out0;
assign v$MUX3_2997_out0 = v$2_2917_out0 ? v$C12_2310_out0 : v$MUX4_725_out0;
assign v$1_3427_out0 = v$G61_3941_out0;
assign v$_5167_out0 = v$MUX7_4758_out0[5:0];
assign v$_5167_out1 = v$MUX7_4758_out0[21:16];
assign v$_361_out0 = { v$2_2917_out0,v$1_3427_out0 };
assign v$MUX2_1039_out0 = v$1_3427_out0 ? v$C13_1292_out0 : v$MUX3_2997_out0;
assign v$X15_2619_out0 = v$_5167_out0;
assign v$_3926_out0 = { v$_5167_out1,v$C2_3735_out0 };
assign v$0_4363_out0 = v$G64_2688_out0;
assign v$SERIESCONNECT_4605_out0 = v$G65_130_out0;
assign v$_483_out0 = { v$0_4363_out0,v$1_3427_out0 };
assign v$_1001_out0 = { v$_20_out0,v$_361_out0 };
assign v$MUX1_2932_out0 = v$0_4363_out0 ? v$C14_2740_out0 : v$MUX2_1039_out0;
assign v$SERIESCONNECT_3100_out0 = v$SERIESCONNECT_4605_out0;
assign v$MUX12_4718_out0 = v$6_1563_out0 ? v$_3926_out0 : v$MUX7_4758_out0;
assign v$SHIFTNUMBER_336_out0 = v$MUX1_2932_out0;
assign v$_1178_out0 = { v$_483_out0,v$2_2917_out0 };
assign v$G41_1467_out0 = v$G45_2792_out0 && v$SERIESCONNECT_3100_out0;
assign v$G43_2434_out0 = v$SEL14_1154_out0 && v$SERIESCONNECT_3100_out0;
assign v$_3605_out0 = { v$_1001_out0,v$0_4363_out0 };
assign v$_4095_out0 = v$MUX12_4718_out0[6:0];
assign v$_4095_out1 = v$MUX12_4718_out0[21:15];
assign v$_2423_out0 = { v$_2315_out0,v$_3605_out0 };
assign v$NOTUSE_2579_out0 = v$SHIFTNUMBER_336_out0;
assign v$X22_2650_out0 = v$_4095_out0;
assign v$G48_2726_out0 = v$G46_560_out0 && v$G41_1467_out0;
assign v$G44_3210_out0 = v$SEL13_3456_out0 && v$G41_1467_out0;
assign v$_3621_out0 = { v$_1178_out0,v$3_4626_out0 };
assign v$_3708_out0 = { v$_4095_out1,v$C9_4326_out0 };
assign v$7_4952_out0 = v$G43_2434_out0;
assign v$G49_3413_out0 = v$SEL16_4039_out0 && v$G48_2726_out0;
assign v$6_3496_out0 = v$G44_3210_out0;
assign v$MUX4_3839_out0 = v$7_1310_out0 ? v$_3708_out0 : v$MUX12_4718_out0;
assign v$G47_4374_out0 = v$G51_3596_out0 && v$G48_2726_out0;
assign v$_4449_out0 = { v$_3621_out0,v$4_1200_out0 };
assign v$OUTPUTSHIFT_5149_out0 = v$_2423_out0;
assign v$G50_247_out0 = v$SEL15_468_out0 && v$G47_4374_out0;
assign v$_747_out0 = v$MUX4_3839_out0[7:0];
assign v$_747_out1 = v$MUX4_3839_out0[21:14];
assign v$_1209_out0 = { v$_4449_out0,v$5_4219_out0 };
assign v$NOTUSE1_1564_out0 = v$OUTPUTSHIFT_5149_out0;
assign v$G54_2009_out0 = v$G52_302_out0 && v$G47_4374_out0;
assign v$5_4220_out0 = v$G49_3413_out0;
assign v$_157_out0 = { v$_747_out1,v$C5_4673_out0 };
assign v$_159_out0 = { v$_1209_out0,v$6_3495_out0 };
assign v$4_1201_out0 = v$G50_247_out0;
assign v$G53_2296_out0 = v$G57_4884_out0 && v$G54_2009_out0;
assign v$G55_3408_out0 = v$SEL18_25_out0 && v$G54_2009_out0;
assign v$X4_4257_out0 = v$_747_out0;
assign v$_4789_out0 = { v$6_3496_out0,v$5_4220_out0 };
assign v$MUX5_156_out0 = v$8_1684_out0 ? v$_157_out0 : v$MUX4_3839_out0;
assign v$G56_2855_out0 = v$SEL17_3945_out0 && v$G53_2296_out0;
assign v$_3121_out0 = { v$7_4952_out0,v$_4789_out0 };
assign v$_3358_out0 = { v$_159_out0,v$7_4951_out0 };
assign v$3_4627_out0 = v$G55_3408_out0;
assign v$G60_5427_out0 = v$G58_4584_out0 && v$G53_2296_out0;
assign v$_21_out0 = { v$4_1201_out0,v$3_4627_out0 };
assign v$_106_out0 = { v$_3358_out0,v$8_1972_out0 };
assign v$G63_822_out0 = v$G62_4942_out0 && v$G60_5427_out0;
assign v$2_2918_out0 = v$G56_2855_out0;
assign v$_3003_out0 = v$MUX5_156_out0[8:0];
assign v$_3003_out1 = v$MUX5_156_out0[21:13];
assign v$G61_3942_out0 = v$SEL20_2271_out0 && v$G60_5427_out0;
assign v$_1290_out0 = { v$_106_out0,v$9_2615_out0 };
assign v$G64_2689_out0 = v$G63_822_out0 && v$SEL21_2092_out0;
assign v$_2838_out0 = { v$_3003_out1,v$C12_4493_out0 };
assign v$1_3428_out0 = v$G61_3942_out0;
assign v$X20_4003_out0 = v$_3003_out0;
assign v$_362_out0 = { v$2_2918_out0,v$1_3428_out0 };
assign v$_933_out0 = { v$_1290_out0,v$10_548_out0 };
assign v$MUX6_1531_out0 = v$9_3255_out0 ? v$_2838_out0 : v$MUX5_156_out0;
assign v$0_4364_out0 = v$G64_2689_out0;
assign v$_484_out0 = { v$0_4364_out0,v$1_3428_out0 };
assign v$_1002_out0 = { v$_21_out0,v$_362_out0 };
assign v$_4578_out0 = v$MUX6_1531_out0[9:0];
assign v$_4578_out1 = v$MUX6_1531_out0[21:12];
assign v$_5398_out0 = { v$_933_out0,v$11_4305_out0 };
assign v$_600_out0 = { v$_5398_out0,v$12_5202_out0 };
assign v$_1179_out0 = { v$_484_out0,v$2_2918_out0 };
assign v$X10_2362_out0 = v$_4578_out0;
assign v$_3606_out0 = { v$_1002_out0,v$0_4364_out0 };
assign v$_5250_out0 = { v$_4578_out1,v$C7_311_out0 };
assign v$MUX3_1699_out0 = v$10_170_out0 ? v$_5250_out0 : v$MUX6_1531_out0;
assign v$OUTPUT_1819_out0 = v$_600_out0;
assign v$_2424_out0 = { v$_3121_out0,v$_3606_out0 };
assign v$_3622_out0 = { v$_1179_out0,v$3_4627_out0 };
assign v$_3067_out0 = v$MUX3_1699_out0[10:0];
assign v$_3067_out1 = v$MUX3_1699_out0[21:11];
assign v$_4450_out0 = { v$_3622_out0,v$4_1201_out0 };
assign v$OUTPUTSHIFT_5150_out0 = v$_2424_out0;
assign v$_1210_out0 = { v$_4450_out0,v$5_4220_out0 };
assign v$_2456_out0 = { v$_3067_out1,v$C11_1736_out0 };
assign v$NOTUSE2_3657_out0 = v$OUTPUTSHIFT_5150_out0;
assign v$X16_4534_out0 = v$_3067_out0;
assign v$_160_out0 = { v$_1210_out0,v$6_3496_out0 };
assign v$MUX10_1398_out0 = v$TOOSMALL_4217_out0 ? v$_2456_out0 : v$MUX3_1699_out0;
assign v$OUT1_1685_out0 = v$MUX10_1398_out0;
assign v$_3359_out0 = { v$_160_out0,v$7_4952_out0 };
assign v$OUTPUT_1820_out0 = v$_3359_out0;
assign v$_728_out0 = { v$OUTPUT_1820_out0,v$OUTPUT_1819_out0 };
assign v$OUTPUT_5043_out0 = v$_728_out0;
assign v$SEL8_352_out0 = v$OUTPUT_5043_out0[8:8];
assign v$SEL9_507_out0 = v$OUTPUT_5043_out0[0:0];
assign v$SEL16_1170_out0 = v$OUTPUT_5043_out0[15:15];
assign v$SEL22_1249_out0 = v$OUTPUT_5043_out0[14:14];
assign v$SEL5_1923_out0 = v$OUTPUT_5043_out0[2:2];
assign v$SEL6_2071_out0 = v$OUTPUT_5043_out0[12:12];
assign v$SEL1_2413_out0 = v$OUTPUT_5043_out0[5:5];
assign v$SEL2_2432_out0 = v$OUTPUT_5043_out0[3:3];
assign v$SEL11_2553_out0 = v$OUTPUT_5043_out0[10:10];
assign v$SEL7_2971_out0 = v$OUTPUT_5043_out0[11:11];
assign v$SEL26_3130_out0 = v$OUTPUT_5043_out0[19:19];
assign v$SEL19_3244_out0 = v$OUTPUT_5043_out0[16:16];
assign v$SEL10_3410_out0 = v$OUTPUT_5043_out0[1:1];
assign v$SEL18_3444_out0 = v$OUTPUT_5043_out0[18:18];
assign v$SEL12_3895_out0 = v$OUTPUT_5043_out0[9:9];
assign v$SEL13_3911_out0 = v$OUTPUT_5043_out0[4:4];
assign v$SEL25_4211_out0 = v$OUTPUT_5043_out0[20:20];
assign v$SEL3_4770_out0 = v$OUTPUT_5043_out0[7:7];
assign v$SEL24_4859_out0 = v$OUTPUT_5043_out0[17:17];
assign v$SEL15_4950_out0 = v$OUTPUT_5043_out0[13:13];
assign v$SEL4_5071_out0 = v$OUTPUT_5043_out0[6:6];
assign v$4_92_out0 = v$SEL13_3911_out0;
assign v$18_146_out0 = v$SEL18_3444_out0;
assign v$15_287_out0 = v$SEL16_1170_out0;
assign v$17_364_out0 = v$SEL24_4859_out0;
assign v$19_506_out0 = v$SEL26_3130_out0;
assign v$6_577_out0 = v$SEL4_5071_out0;
assign v$5_720_out0 = v$SEL1_2413_out0;
assign v$3_875_out0 = v$SEL2_2432_out0;
assign v$7_1058_out0 = v$SEL3_4770_out0;
assign v$13_1171_out0 = v$SEL15_4950_out0;
assign v$2_1456_out0 = v$SEL5_1923_out0;
assign v$0_1730_out0 = v$SEL9_507_out0;
assign v$10_1774_out0 = v$SEL11_2553_out0;
assign v$16_1807_out0 = v$SEL19_3244_out0;
assign v$1_1838_out0 = v$SEL10_3410_out0;
assign v$14_2190_out0 = v$SEL22_1249_out0;
assign v$9_2870_out0 = v$SEL12_3895_out0;
assign v$8_3011_out0 = v$SEL8_352_out0;
assign v$12_3049_out0 = v$SEL6_2071_out0;
assign v$20_3698_out0 = v$SEL25_4211_out0;
assign v$11_5022_out0 = v$SEL7_2971_out0;
assign v$MUX4_5413_out0 = v$20_3698_out0 ? v$C10_3628_out0 : v$C10_3628_out0;
assign v$MUX12_4936_out0 = v$19_506_out0 ? v$C13_5266_out0 : v$MUX4_5413_out0;
assign v$MUX13_1767_out0 = v$18_146_out0 ? v$C1_4327_out0 : v$MUX12_4936_out0;
assign v$MUX2_5303_out0 = v$17_364_out0 ? v$C11_3973_out0 : v$MUX13_1767_out0;
assign v$MUX7_685_out0 = v$16_1807_out0 ? v$C12_1322_out0 : v$MUX2_5303_out0;
assign v$MUX8_4023_out0 = v$15_287_out0 ? v$C3_1385_out0 : v$MUX7_685_out0;
assign v$MUX11_5024_out0 = v$14_2190_out0 ? v$C6_34_out0 : v$MUX8_4023_out0;
assign v$MUX6_3257_out0 = v$13_1171_out0 ? v$C8_3052_out0 : v$MUX11_5024_out0;
assign v$MUX1_493_out0 = v$12_3049_out0 ? v$C4_3256_out0 : v$MUX6_3257_out0;
assign v$MUX22_5423_out0 = v$11_5022_out0 ? v$C19_5406_out0 : v$MUX1_493_out0;
assign v$MUX19_2194_out0 = v$10_1774_out0 ? v$C22_372_out0 : v$MUX22_5423_out0;
assign v$MUX16_4015_out0 = v$9_2870_out0 ? v$C21_5199_out0 : v$MUX19_2194_out0;
assign v$MUX21_3934_out0 = v$8_3011_out0 ? v$C20_1438_out0 : v$MUX16_4015_out0;
assign v$MUX15_1450_out0 = v$7_1058_out0 ? v$C15_2147_out0 : v$MUX21_3934_out0;
assign v$MUX18_5418_out0 = v$6_577_out0 ? v$C16_427_out0 : v$MUX15_1450_out0;
assign v$MUX20_4105_out0 = v$5_720_out0 ? v$C14_576_out0 : v$MUX18_5418_out0;
assign v$MUX17_3354_out0 = v$4_92_out0 ? v$C17_1139_out0 : v$MUX20_4105_out0;
assign v$MUX14_3139_out0 = v$3_875_out0 ? v$C18_3898_out0 : v$MUX17_3354_out0;
assign v$MUX31_1588_out0 = v$2_1456_out0 ? v$C28_1010_out0 : v$MUX14_3139_out0;
assign v$MUX28_810_out0 = v$1_1838_out0 ? v$C31_3551_out0 : v$MUX31_1588_out0;
assign v$MUX25_5182_out0 = v$0_1730_out0 ? v$C30_4304_out0 : v$MUX28_810_out0;
assign v$SHIFTNUMBER_3013_out0 = v$MUX25_5182_out0;
assign v$SHIFTNUMBER_5176_out0 = v$SHIFTNUMBER_3013_out0;
assign v$SHIFTNUMBER_3952_out0 = v$SHIFTNUMBER_5176_out0;
assign v$_2649_out0 = { v$SHIFTNUMBER_3952_out0,v$C31_1111_out0 };
assign v$_3086_out0 = { v$SHIFTNUMBER_3952_out0,v$C18_1515_out0 };
assign v$XOR1_3485_out0 = v$_3086_out0 ^ v$C15_3896_out0;
assign {v$A1_2125_out1,v$A1_2125_out0 } = v$_2023_out0 + v$XOR1_3485_out0 + v$C14_4932_out0;
assign v$_862_out0 = v$A1_2125_out0[6:0];
assign v$_862_out1 = v$A1_2125_out0[7:1];
assign v$COUT_1150_out0 = v$A1_2125_out1;
assign v$EQ15_2420_out0 = v$A1_2125_out0 == 8'h0;
assign v$DIFFERENCE7_132_out0 = v$_862_out0;
assign v$EQ16_329_out0 = v$_862_out1 == 1'h0;
assign v$EQUAL_5338_out0 = v$EQ15_2420_out0;
assign v$SEL4_464_out0 = v$DIFFERENCE7_132_out0[5:5];
assign v$EXPOBIGGER_2482_out0 = v$EQ16_329_out0;
assign v$SEL3_3088_out0 = v$DIFFERENCE7_132_out0[6:6];
assign v$SEL2_3828_out0 = v$DIFFERENCE7_132_out0[4:0];
assign v$MUX14_141_out0 = v$EXPOBIGGER_2482_out0 ? v$_2649_out0 : v$EXPONENT_5089_out0;
assign v$G1_2937_out0 = ! v$SEL3_3088_out0;
assign v$EQ26_4856_out0 = v$SEL2_3828_out0 == 5'h1f;
assign v$DIFFERENCE_5352_out0 = v$SEL2_3828_out0;
assign v$MUX16_907_out0 = v$EQUAL_5338_out0 ? v$C17_5302_out0 : v$DIFFERENCE_5352_out0;
assign v$SHIFT_3099_out0 = v$MUX14_141_out0;
assign v$G3_3808_out0 = v$SEL4_464_out0 || v$EQ26_4856_out0;
assign v$EQ17_35_out0 = v$SHIFT_3099_out0 == 7'h12;
assign v$EQ7_379_out0 = v$SHIFT_3099_out0 == 7'h5;
assign v$G2_704_out0 = v$G1_2937_out0 && v$G3_3808_out0;
assign v$EQ11_707_out0 = v$SHIFT_3099_out0 == 7'ha;
assign v$EQ25_1034_out0 = v$SHIFT_3099_out0 == 7'h10;
assign v$EQ20_1460_out0 = v$SHIFT_3099_out0 == 7'hf;
assign v$EQ24_1543_out0 = v$SHIFT_3099_out0 == 7'h14;
assign v$EQ5_1712_out0 = v$SHIFT_3099_out0 == 7'h4;
assign v$EQ22_1837_out0 = v$SHIFT_3099_out0 == 7'he;
assign v$EQ1_1858_out0 = v$SHIFT_3099_out0 == 7'h0;
assign v$EQ12_2481_out0 = v$SHIFT_3099_out0 == 7'hb;
assign v$EQ9_2487_out0 = v$SHIFT_3099_out0 == 7'h9;
assign v$EQ18_3008_out0 = v$SHIFT_3099_out0 == 7'h11;
assign v$EQ3_3281_out0 = v$SHIFT_3099_out0 == 7'h2;
assign v$EQ6_3801_out0 = v$SHIFT_3099_out0 == 7'h6;
assign v$EQ2_4098_out0 = v$SHIFT_3099_out0 == 7'h1;
assign v$EQ21_4249_out0 = v$SHIFT_3099_out0 == 7'h13;
assign v$EQ10_4417_out0 = v$SHIFT_3099_out0 == 7'h8;
assign v$EQ19_4433_out0 = v$SHIFT_3099_out0 == 7'hd;
assign v$EQ8_5195_out0 = v$SHIFT_3099_out0 == 7'h7;
assign v$MUX15_5222_out0 = v$EXPOBIGGER_2482_out0 ? v$MUX16_907_out0 : v$C16_205_out0;
assign v$EQ13_5289_out0 = v$SHIFT_3099_out0 == 7'hc;
assign v$EQ4_5388_out0 = v$SHIFT_3099_out0 == 7'h3;
assign v$15_2_out0 = v$EQ20_1460_out0;
assign v$19_240_out0 = v$EQ21_4249_out0;
assign v$6_324_out0 = v$EQ6_3801_out0;
assign v$8_401_out0 = v$EQ10_4417_out0;
assign v$9_784_out0 = v$EQ9_2487_out0;
assign v$14_1168_out0 = v$EQ22_1837_out0;
assign v$11_1205_out0 = v$EQ12_2481_out0;
assign v$2_1286_out0 = v$EQ3_3281_out0;
assign v$NEWEXPONENT_1710_out0 = v$MUX15_5222_out0;
assign v$7_1771_out0 = v$EQ8_5195_out0;
assign v$4_2368_out0 = v$EQ5_1712_out0;
assign v$16_2631_out0 = v$EQ25_1034_out0;
assign v$12_2738_out0 = v$EQ13_5289_out0;
assign v$OVERFLOW_2773_out0 = v$G2_704_out0;
assign v$13_3103_out0 = v$EQ19_4433_out0;
assign v$20_3805_out0 = v$EQ24_1543_out0;
assign v$17_4021_out0 = v$EQ18_3008_out0;
assign v$18_4283_out0 = v$EQ17_35_out0;
assign v$10_4288_out0 = v$EQ11_707_out0;
assign v$0_4489_out0 = v$EQ1_1858_out0;
assign v$5_4614_out0 = v$EQ7_379_out0;
assign v$1_5101_out0 = v$EQ2_4098_out0;
assign v$3_5238_out0 = v$EQ4_5388_out0;
assign v$MUX1_533_out0 = v$1_5101_out0 ? v$_416_out0 : v$_2865_out0;
assign v$NEWEXPO0001_1724_out0 = v$NEWEXPONENT_1710_out0;
assign v$OVERFLOW0_5258_out0 = v$OVERFLOW_2773_out0;
assign v$MUX2_37_out0 = v$MULTISHIFT_2679_out0 ? v$NEWEXPO0001_1724_out0 : v$NEWEXPO1011_4381_out0;
assign v$MUX6_572_out0 = v$MULTISHIFT_2679_out0 ? v$OVERFLOW0_5258_out0 : v$OVERFLOW1_4085_out0;
assign v$_3525_out0 = v$MUX1_533_out0[18:0];
assign v$_3525_out1 = v$MUX1_533_out0[20:2];
assign v$G4_597_out0 = v$MUX6_572_out0 || v$INFINITY_1025_out0;
assign v$X1_816_out0 = v$_3525_out1;
assign v$MUX1_3829_out0 = v$NEGATIVEMODE_394_out0 ? v$C1_2206_out0 : v$MUX2_37_out0;
assign v$_5424_out0 = { v$C3_3893_out0,v$_3525_out0 };
assign v$EXCEPTION_1020_out0 = v$G4_597_out0;
assign v$EXPO0IFNEG_1045_out0 = v$MUX1_3829_out0;
assign v$EXCEPTION_1689_out0 = v$G4_597_out0;
assign v$MUX2_3635_out0 = v$2_1286_out0 ? v$_5424_out0 : v$MUX1_533_out0;
assign v$G9_567_out0 = v$EXCEPTION_5275_out0 || v$EXCEPTION_1689_out0;
assign v$_3618_out0 = v$MUX2_3635_out0[17:0];
assign v$_3618_out1 = v$MUX2_3635_out0[20:3];
assign v$MUX5_3998_out0 = v$EXCEPTION_1020_out0 ? v$C2_2234_out0 : v$EXPO0IFNEG_1045_out0;
assign v$_33_out0 = { v$C4_627_out0,v$_3618_out0 };
assign v$X2_531_out0 = v$_3618_out1;
assign v$EXCEPTION_1402_out0 = v$G9_567_out0;
assign v$NEWEXPO_5072_out0 = v$MUX5_3998_out0;
assign v$EXCEPTION_321_out0 = v$EXCEPTION_1402_out0;
assign v$MUX3_5301_out0 = v$3_5238_out0 ? v$_33_out0 : v$MUX2_3635_out0;
assign v$EXCEPTION_1252_out0 = v$EXCEPTION_321_out0;
assign v$_3740_out0 = v$MUX3_5301_out0[16:0];
assign v$_3740_out1 = v$MUX3_5301_out0[20:4];
assign v$X3_1541_out0 = v$_3740_out1;
assign v$_5389_out0 = { v$C5_4214_out0,v$_3740_out0 };
assign v$MUX4_3788_out0 = v$4_2368_out0 ? v$_5389_out0 : v$MUX3_5301_out0;
assign v$_2089_out0 = v$MUX4_3788_out0[15:0];
assign v$_2089_out1 = v$MUX4_3788_out0[20:5];
assign v$X5_134_out0 = v$_2089_out1;
assign v$_3261_out0 = { v$C6_3198_out0,v$_2089_out0 };
assign v$MUX5_3531_out0 = v$5_4614_out0 ? v$_3261_out0 : v$MUX4_3788_out0;
assign v$_4372_out0 = v$MUX5_3531_out0[14:0];
assign v$_4372_out1 = v$MUX5_3531_out0[20:6];
assign v$_2131_out0 = { v$C7_228_out0,v$_4372_out0 };
assign v$X4_3285_out0 = v$_4372_out1;
assign v$MUX6_5312_out0 = v$6_324_out0 ? v$_2131_out0 : v$MUX5_3531_out0;
assign v$_3090_out0 = v$MUX6_5312_out0[13:0];
assign v$_3090_out1 = v$MUX6_5312_out0[20:7];
assign v$_0_out0 = { v$C8_4082_out0,v$_3090_out0 };
assign v$X7_4476_out0 = v$_3090_out1;
assign v$MUX8_1156_out0 = v$7_1771_out0 ? v$_0_out0 : v$MUX6_5312_out0;
assign v$_1278_out0 = v$MUX8_1156_out0[12:0];
assign v$_1278_out1 = v$MUX8_1156_out0[20:8];
assign v$X6_230_out0 = v$_1278_out1;
assign v$_3128_out0 = { v$C9_758_out0,v$_1278_out0 };
assign v$MUX7_1475_out0 = v$8_401_out0 ? v$_3128_out0 : v$MUX8_1156_out0;
assign v$_2309_out0 = v$MUX7_1475_out0[11:0];
assign v$_2309_out1 = v$MUX7_1475_out0[20:9];
assign v$X8_4348_out0 = v$_2309_out1;
assign v$_4773_out0 = { v$C10_5296_out0,v$_2309_out0 };
assign v$MUX9_2441_out0 = v$9_784_out0 ? v$_4773_out0 : v$MUX7_1475_out0;
assign v$_1145_out0 = v$MUX9_2441_out0[10:0];
assign v$_1145_out1 = v$MUX9_2441_out0[20:10];
assign v$X17_1251_out0 = v$_1145_out1;
assign v$_2422_out0 = { v$C12_3681_out0,v$_1145_out0 };
assign v$MUX11_990_out0 = v$10_4288_out0 ? v$_2422_out0 : v$MUX9_2441_out0;
assign v$_1361_out0 = v$MUX11_990_out0[9:0];
assign v$_1361_out1 = v$MUX11_990_out0[20:11];
assign v$_1241_out0 = { v$C11_4416_out0,v$_1361_out0 };
assign v$X13_3686_out0 = v$_1361_out1;
assign v$MUX12_4386_out0 = v$11_1205_out0 ? v$_1241_out0 : v$MUX11_990_out0;
assign v$_1016_out0 = v$MUX12_4386_out0[8:0];
assign v$_1016_out1 = v$MUX12_4386_out0[20:12];
assign v$X16_4303_out0 = v$_1016_out1;
assign v$_5248_out0 = { v$C13_325_out0,v$_1016_out0 };
assign v$MUX13_300_out0 = v$12_2738_out0 ? v$_5248_out0 : v$MUX12_4386_out0;
assign v$_1387_out0 = v$MUX13_300_out0[7:0];
assign v$_1387_out1 = v$MUX13_300_out0[20:13];
assign v$X21_241_out0 = v$_1387_out1;
assign v$_588_out0 = { v$C21_4143_out0,v$_1387_out0 };
assign v$MUX18_2756_out0 = v$13_3103_out0 ? v$_588_out0 : v$MUX13_300_out0;
assign v$_3556_out0 = v$MUX18_2756_out0[6:0];
assign v$_3556_out1 = v$MUX18_2756_out0[20:14];
assign v$X24_2269_out0 = v$_3556_out1;
assign v$_5245_out0 = { v$C28_4909_out0,v$_3556_out0 };
assign v$MUX24_3282_out0 = v$14_1168_out0 ? v$_5245_out0 : v$MUX18_2756_out0;
assign v$_1688_out0 = v$MUX24_3282_out0[5:0];
assign v$_1688_out1 = v$MUX24_3282_out0[20:15];
assign v$X22_626_out0 = v$_1688_out1;
assign v$_4446_out0 = { v$C24_4122_out0,v$_1688_out0 };
assign v$MUX27_2678_out0 = v$15_2_out0 ? v$_4446_out0 : v$MUX24_3282_out0;
assign v$_4691_out0 = v$MUX27_2678_out0[4:0];
assign v$_4691_out1 = v$MUX27_2678_out0[20:16];
assign v$X27_3311_out0 = v$_4691_out1;
assign v$_5032_out0 = { v$C30_3636_out0,v$_4691_out0 };
assign v$MUX25_1038_out0 = v$16_2631_out0 ? v$_5032_out0 : v$MUX27_2678_out0;
assign v$_4475_out0 = v$MUX25_1038_out0[3:0];
assign v$_4475_out1 = v$MUX25_1038_out0[20:17];
assign v$_635_out0 = { v$C26_791_out0,v$_4475_out0 };
assign v$X18_2941_out0 = v$_4475_out1;
assign v$MUX23_3043_out0 = v$17_4021_out0 ? v$_635_out0 : v$MUX25_1038_out0;
assign v$_3677_out0 = v$MUX23_3043_out0[2:0];
assign v$_3677_out1 = v$MUX23_3043_out0[20:18];
assign v$_1906_out0 = { v$C22_4676_out0,v$_3677_out0 };
assign v$X31_4020_out0 = v$_3677_out1;
assign v$MUX28_5060_out0 = v$18_4283_out0 ? v$_1906_out0 : v$MUX23_3043_out0;
assign v$_4862_out0 = v$MUX28_5060_out0[1:0];
assign v$_4862_out1 = v$MUX28_5060_out0[20:19];
assign v$X38_1004_out0 = v$_4862_out1;
assign v$_5220_out0 = { v$C29_4076_out0,v$_4862_out0 };
assign v$MUX20_5281_out0 = v$19_240_out0 ? v$_5220_out0 : v$MUX28_5060_out0;
assign v$_4931_out0 = v$MUX20_5281_out0[0:0];
assign v$_4931_out1 = v$MUX20_5281_out0[20:20];
assign v$X20_2699_out0 = v$_4931_out1;
assign v$_4415_out0 = { v$C25_3012_out0,v$_4931_out0 };
assign v$MUX21_762_out0 = v$20_3805_out0 ? v$_4415_out0 : v$MUX20_5281_out0;
assign v$_2772_out0 = { v$MUX21_762_out0,v$C32_2090_out0 };
assign v$OUT_3656_out0 = v$_2772_out0;
assign v$NEWFRAC0001_4382_out0 = v$OUT_3656_out0;
assign v$MUX3_4210_out0 = v$MULTISHIFT_2679_out0 ? v$NEWFRAC0001_4382_out0 : v$NEWFRAC1011_2046_out0;
assign v$MUX4_48_out0 = v$NEGATIVEMODE_394_out0 ? v$OUT1_1685_out0 : v$MUX3_4210_out0;
assign v$_691_out0 = v$MUX4_48_out0[9:0];
assign v$_691_out1 = v$MUX4_48_out0[21:12];
assign v$ROUNDEDBITS_4566_out0 = v$_691_out0;
assign v$_4938_out0 = v$_691_out1[9:0];
assign v$_4938_out1 = v$_691_out1[11:2];
assign v$MUX7_1172_out0 = v$EXCEPTION_1020_out0 ? v$C4_268_out0 : v$_4938_out0;
assign v$INT_4565_out0 = v$_4938_out1;
assign v$NEWFRAC_3836_out0 = v$MUX7_1172_out0;
assign v$_328_out0 = { v$NEWFRAC_3836_out0,v$NEWEXPO_5072_out0 };
assign v$_5152_out0 = { v$_328_out0,v$SGN_3620_out0 };
assign v$MUX1_3947_out0 = v$MULT_991_out0 ? v$_5152_out0 : v$fpmerge_5196_out0;
assign v$FPOUT_4479_out0 = v$MUX1_3947_out0;
assign v$MUX2_5187_out0 = v$CYC2_1461_out0 ? v$FPOUT_4479_out0 : v$WDATA_4407_out0;


endmodule
