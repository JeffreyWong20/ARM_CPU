
module main (
	clk,
	v$READVALID_17_out0,
	v$WRITECOMPLETE_55_out0,
	v$INTERRUPT_418_out0,
	v$PCORROM_461_out0,
	v$PRIORITY_333_out0,
	v$R3_251_out0,
	v$R2_370_out0,
	v$R0_525_out0,
	v$R1_691_out0,
	v$PROGRAMADDRESS_616_out0);
input clk;
input  [15:0] v$PCORROM_461_out0;
input v$INTERRUPT_418_out0;
input v$READVALID_17_out0;
input v$WRITECOMPLETE_55_out0;
output  [11:0] v$PROGRAMADDRESS_616_out0;
output  [15:0] v$R0_525_out0;
output  [15:0] v$R1_691_out0;
output  [15:0] v$R2_370_out0;
output  [15:0] v$R3_251_out0;
output v$PRIORITY_333_out0;
reg  [11:0] v$REG1_43_out0 = 12'h0;
reg  [11:0] v$REG2_86_out0 = 12'h0;
reg  [15:0] v$REG0_622_out0 = 16'h0;
reg  [15:0] v$REG1_164_out0 = 16'h0;
reg  [15:0] v$REG1_339_out0 = 16'h0;
reg  [15:0] v$REG1_434_out0 = 16'h0;
reg  [15:0] v$REG1_485_out0 = 16'h0;
reg  [15:0] v$REG2_355_out0 = 16'h0;
reg  [15:0] v$REG2_665_out0 = 16'h0;
reg  [15:0] v$REG3_263_out0 = 16'h0;
reg  [15:0] v$REG3_383_out0 = 16'h0;
reg  [15:0] v$REG4_215_out0 = 16'h0;
reg  [15:0] v$REG4_660_out0 = 16'h0;
reg  [15:0] v$REG5_394_out0 = 16'h0;
reg v$FF1_14_out0 = 1'b0;
reg v$FF1_186_out0 = 1'b0;
reg v$FF1_192_out0 = 1'b0;
reg v$FF1_248_out0 = 1'b0;
reg v$FF1_386_out0 = 1'b0;
reg v$FF1_564_out0 = 1'b0;
reg v$FF2_325_out0 = 1'b0;
reg v$FF2_437_out0 = 1'b0;
reg v$FF2_570_out0 = 1'b0;
reg v$FF2_601_out0 = 1'b0;
reg v$FF3_606_out0 = 1'b0;
reg v$FF4_416_out0 = 1'b0;
reg v$REG2_235_out0 = 1'b0;
reg v$REG3_65_out0 = 1'b0;
wire  [10:0] v$C1_141_out0;
wire  [10:0] v$_387_out1;
wire  [10:0] v$_698_out1;
wire  [11:0] v$A1_369_out0;
wire  [11:0] v$C1_209_out0;
wire  [11:0] v$C1_245_out0;
wire  [11:0] v$C4_406_out0;
wire  [11:0] v$IR110_675_out0;
wire  [11:0] v$IR12_436_out0;
wire  [11:0] v$MUX1_531_out0;
wire  [11:0] v$MUX2_87_out0;
wire  [11:0] v$MUX4_89_out0;
wire  [11:0] v$MUX5_366_out0;
wire  [11:0] v$MUX6_456_out0;
wire  [11:0] v$MUX7_592_out0;
wire  [11:0] v$N_681_out0;
wire  [11:0] v$PC1_115_out0;
wire  [11:0] v$PC_590_out0;
wire  [11:0] v$RAMADDRMUX_173_out0;
wire  [11:0] v$RAMADDRMUX_505_out0;
wire  [11:0] v$RAMADDRMUX_723_out0;
wire  [11:0] v$RAMADDRMUX_72_out0;
wire  [11:0] v$STOREDPC_415_out0;
wire  [11:0] v$STOREDPC_718_out0;
wire  [11:0] v$_202_out1;
wire  [11:0] v$_358_out1;
wire  [11:0] v$_411_out1;
wire  [11:0] v$_444_out0;
wire  [11:0] v$_454_out0;
wire  [11:0] v$_614_out0;
wire  [12:0] v$_150_out1;
wire  [12:0] v$_272_out1;
wire  [13:0] v$_129_out0;
wire  [13:0] v$_1_out1;
wire  [13:0] v$_207_out1;
wire  [13:0] v$_602_out1;
wire  [14:0] v$_25_out1;
wire  [14:0] v$_287_out0;
wire  [14:0] v$_470_out0;
wire  [14:0] v$_501_out1;
wire  [14:0] v$_672_out1;
wire  [14:0] v$_99_out1;
wire  [15:0] v$1TO4_487_out0;
wire  [15:0] v$A1_135_out0;
wire  [15:0] v$A1_38_out0;
wire  [15:0] v$ALUOUT_174_out0;
wire  [15:0] v$ALUOUT_214_out0;
wire  [15:0] v$ALUOUT_477_out0;
wire  [15:0] v$ALUOUT_506_out0;
wire  [15:0] v$ALUOUT_61_out0;
wire  [15:0] v$ALUOUT_721_out0;
wire  [15:0] v$ANDOUT_460_out0;
wire  [15:0] v$ASR_22_out0;
wire  [15:0] v$ASR_377_out0;
wire  [15:0] v$ASR_76_out0;
wire  [15:0] v$ASR_93_out0;
wire  [15:0] v$A_656_out0;
wire  [15:0] v$B_558_out0;
wire  [15:0] v$C1_97_out0;
wire  [15:0] v$C2_743_out0;
wire  [15:0] v$C3_179_out0;
wire  [15:0] v$C4_46_out0;
wire  [15:0] v$DIN3_518_out0;
wire  [15:0] v$DOUT1_98_out0;
wire  [15:0] v$DOUT2_117_out0;
wire  [15:0] v$EA_341_out0;
wire  [15:0] v$IN_120_out0;
wire  [15:0] v$IN_222_out0;
wire  [15:0] v$IN_307_out0;
wire  [15:0] v$IN_310_out0;
wire  [15:0] v$IN_384_out0;
wire  [15:0] v$IN_412_out0;
wire  [15:0] v$IN_41_out0;
wire  [15:0] v$IN_619_out0;
wire  [15:0] v$IN_626_out0;
wire  [15:0] v$IN_667_out0;
wire  [15:0] v$IN_673_out0;
wire  [15:0] v$IR16_716_out0;
wire  [15:0] v$IR_27_out0;
wire  [15:0] v$IR_297_out0;
wire  [15:0] v$IR_330_out0;
wire  [15:0] v$IR_526_out0;
wire  [15:0] v$IR_94_out0;
wire  [15:0] v$LSL_163_out0;
wire  [15:0] v$LSL_250_out0;
wire  [15:0] v$LSL_515_out0;
wire  [15:0] v$LSL_738_out0;
wire  [15:0] v$LSR_268_out0;
wire  [15:0] v$LSR_335_out0;
wire  [15:0] v$LSR_402_out0;
wire  [15:0] v$LSR_677_out0;
wire  [15:0] v$MSL_68_out0;
wire  [15:0] v$MSR_321_out0;
wire  [15:0] v$MUX10_266_out0;
wire  [15:0] v$MUX11_165_out0;
wire  [15:0] v$MUX12_15_out0;
wire  [15:0] v$MUX13_548_out0;
wire  [15:0] v$MUX14_198_out0;
wire  [15:0] v$MUX1_168_out0;
wire  [15:0] v$MUX1_194_out0;
wire  [15:0] v$MUX1_349_out0;
wire  [15:0] v$MUX1_393_out0;
wire  [15:0] v$MUX1_475_out0;
wire  [15:0] v$MUX1_489_out0;
wire  [15:0] v$MUX1_512_out0;
wire  [15:0] v$MUX1_524_out0;
wire  [15:0] v$MUX1_547_out0;
wire  [15:0] v$MUX1_598_out0;
wire  [15:0] v$MUX1_664_out0;
wire  [15:0] v$MUX1_731_out0;
wire  [15:0] v$MUX2_256_out0;
wire  [15:0] v$MUX2_265_out0;
wire  [15:0] v$MUX2_280_out0;
wire  [15:0] v$MUX2_360_out0;
wire  [15:0] v$MUX2_511_out0;
wire  [15:0] v$MUX2_642_out0;
wire  [15:0] v$MUX2_90_out0;
wire  [15:0] v$MUX3_306_out0;
wire  [15:0] v$MUX3_425_out0;
wire  [15:0] v$MUX3_427_out0;
wire  [15:0] v$MUX3_42_out0;
wire  [15:0] v$MUX3_442_out0;
wire  [15:0] v$MUX3_54_out0;
wire  [15:0] v$MUX3_671_out0;
wire  [15:0] v$MUX3_724_out0;
wire  [15:0] v$MUX4_127_out0;
wire  [15:0] v$MUX4_156_out0;
wire  [15:0] v$MUX4_234_out0;
wire  [15:0] v$MUX4_28_out0;
wire  [15:0] v$MUX4_49_out0;
wire  [15:0] v$MUX4_51_out0;
wire  [15:0] v$MUX4_725_out0;
wire  [15:0] v$MUX5_403_out0;
wire  [15:0] v$MUX5_498_out0;
wire  [15:0] v$MUX6_170_out0;
wire  [15:0] v$MUX6_91_out0;
wire  [15:0] v$MUX7_389_out0;
wire  [15:0] v$MUX8_206_out0;
wire  [15:0] v$MUX9_508_out0;
wire  [15:0] v$OP1_176_out0;
wire  [15:0] v$OP1_555_out0;
wire  [15:0] v$OP2_257_out0;
wire  [15:0] v$OP2_348_out0;
wire  [15:0] v$OP2_388_out0;
wire  [15:0] v$OP2_546_out0;
wire  [15:0] v$OUT_128_out0;
wire  [15:0] v$OUT_212_out0;
wire  [15:0] v$OUT_399_out0;
wire  [15:0] v$OUT_624_out0;
wire  [15:0] v$OUT_730_out0;
wire  [15:0] v$R0S_140_out0;
wire  [15:0] v$R0S_148_out0;
wire  [15:0] v$R0TEST_283_out0;
wire  [15:0] v$R0TEST_700_out0;
wire  [15:0] v$R0_106_out0;
wire  [15:0] v$R0_124_out0;
wire  [15:0] v$R0_519_out0;
wire  [15:0] v$R0_571_out0;
wire  [15:0] v$R1S_29_out0;
wire  [15:0] v$R1S_669_out0;
wire  [15:0] v$R1TEST_376_out0;
wire  [15:0] v$R1TEST_551_out0;
wire  [15:0] v$R1_375_out0;
wire  [15:0] v$R1_490_out0;
wire  [15:0] v$R1_561_out0;
wire  [15:0] v$R1_588_out0;
wire  [15:0] v$R2S_161_out0;
wire  [15:0] v$R2S_467_out0;
wire  [15:0] v$R2TEST_152_out0;
wire  [15:0] v$R2TEST_583_out0;
wire  [15:0] v$R2_264_out0;
wire  [15:0] v$R2_391_out0;
wire  [15:0] v$R2_529_out0;
wire  [15:0] v$R2_687_out0;
wire  [15:0] v$R3S_648_out0;
wire  [15:0] v$R3S_650_out0;
wire  [15:0] v$R3TEST_242_out0;
wire  [15:0] v$R3TEST_732_out0;
wire  [15:0] v$R3_232_out0;
wire  [15:0] v$R3_276_out0;
wire  [15:0] v$R3_363_out0;
wire  [15:0] v$R3_693_out0;
wire  [15:0] v$RAMDOUT_254_out0;
wire  [15:0] v$RAMDOUT_337_out0;
wire  [15:0] v$RAMDOUT_356_out0;
wire  [15:0] v$RAMDOUT_367_out0;
wire  [15:0] v$RAMDOUT_639_out0;
wire  [15:0] v$RDOUT_216_out0;
wire  [15:0] v$RDOUT_33_out0;
wire  [15:0] v$RD_260_out0;
wire  [15:0] v$REGDIN_238_out0;
wire  [15:0] v$REGDIN_446_out0;
wire  [15:0] v$RMN_452_out0;
wire  [15:0] v$RMN_95_out0;
wire  [15:0] v$RM_142_out0;
wire  [15:0] v$RM_210_out0;
wire  [15:0] v$RM_284_out0;
wire  [15:0] v$RM_392_out0;
wire  [15:0] v$RM_458_out0;
wire  [15:0] v$RM_620_out0;
wire  [15:0] v$RM_685_out0;
wire  [15:0] v$ROR_118_out0;
wire  [15:0] v$ROR_201_out0;
wire  [15:0] v$ROR_324_out0;
wire  [15:0] v$ROR_353_out0;
wire  [15:0] v$SHIFTIN_300_out0;
wire  [15:0] v$SHIFTOUT_221_out0;
wire  [15:0] v$XOR1_169_out0;
wire  [15:0] v$XOR1_253_out0;
wire  [15:0] v$X_617_out0;
wire  [15:0] v$_108_out0;
wire  [15:0] v$_109_out0;
wire  [15:0] v$_180_out0;
wire  [15:0] v$_20_out0;
wire  [15:0] v$_224_out0;
wire  [15:0] v$_30_out0;
wire  [15:0] v$_320_out0;
wire  [15:0] v$_395_out0;
wire  [15:0] v$_398_out0;
wire  [15:0] v$_408_out0;
wire  [15:0] v$_44_out0;
wire  [15:0] v$_453_out0;
wire  [15:0] v$_457_out0;
wire  [15:0] v$_481_out0;
wire  [15:0] v$_510_out0;
wire  [15:0] v$_566_out0;
wire  [15:0] v$_567_out0;
wire  [15:0] v$_56_out0;
wire  [15:0] v$_69_out0;
wire  [15:0] v$_728_out0;
wire  [15:0] v$_78_out0;
wire  [1:0] v$2_468_out0;
wire  [1:0] v$3_4_out0;
wire  [1:0] v$6_116_out0;
wire  [1:0] v$8_11_out0;
wire  [1:0] v$9_131_out0;
wire  [1:0] v$AD1_742_out0;
wire  [1:0] v$AD2_581_out0;
wire  [1:0] v$AD3_550_out0;
wire  [1:0] v$C1_540_out0;
wire  [1:0] v$D_359_out0;
wire  [1:0] v$D_59_out0;
wire  [1:0] v$D_707_out0;
wire  [1:0] v$MUX1_3_out0;
wire  [1:0] v$MUX2_112_out0;
wire  [1:0] v$M_138_out0;
wire  [1:0] v$M_629_out0;
wire  [1:0] v$Q1_618_out0;
wire  [1:0] v$Q_517_out0;
wire  [1:0] v$Q_729_out0;
wire  [1:0] v$ROR_430_out0;
wire  [1:0] v$SHIFTPREVIOUS_187_out0;
wire  [1:0] v$SHIFT_182_out0;
wire  [1:0] v$SHIFT_271_out0;
wire  [1:0] v$SR_104_out0;
wire  [1:0] v$SR_317_out0;
wire  [1:0] v$SR_414_out0;
wire  [1:0] v$SR_537_out0;
wire  [1:0] v$SR_565_out0;
wire  [1:0] v$SR_659_out0;
wire  [1:0] v$ZERO_439_out0;
wire  [1:0] v$_123_out0;
wire  [1:0] v$_129_out1;
wire  [1:0] v$_196_out0;
wire  [1:0] v$_205_out0;
wire  [1:0] v$_21_out1;
wire  [1:0] v$_318_out0;
wire  [1:0] v$_322_out0;
wire  [1:0] v$_344_out0;
wire  [1:0] v$_350_out1;
wire  [1:0] v$_463_out0;
wire  [1:0] v$_473_out0;
wire  [1:0] v$_480_out0;
wire  [1:0] v$_520_out0;
wire  [1:0] v$_577_out0;
wire  [1:0] v$_579_out0;
wire  [1:0] v$_602_out0;
wire  [1:0] v$_680_out0;
wire  [1:0] v$_746_out0;
wire  [1:0] v$_88_out1;
wire  [2:0] v$1_597_out0;
wire  [2:0] v$NA_474_out0;
wire  [2:0] v$OP_110_out0;
wire  [2:0] v$OP_58_out0;
wire  [2:0] v$_378_out1;
wire  [2:0] v$_654_out1;
wire  [2:0] v$_694_out0;
wire  [2:0] v$_733_out1;
wire  [3:0] v$4_288_out0;
wire  [3:0] v$5_71_out0;
wire  [3:0] v$9_400_out0;
wire  [3:0] v$B_114_out0;
wire  [3:0] v$B_241_out0;
wire  [3:0] v$B_464_out0;
wire  [3:0] v$B_66_out0;
wire  [3:0] v$C1_486_out0;
wire  [3:0] v$NOTUSED_649_out0;
wire  [3:0] v$N_343_out0;
wire  [3:0] v$N_715_out0;
wire  [3:0] v$O_312_out0;
wire  [3:0] v$SEL1_64_out0;
wire  [3:0] v$ZERO_426_out0;
wire  [3:0] v$_155_out1;
wire  [3:0] v$_177_out0;
wire  [3:0] v$_294_out0;
wire  [3:0] v$_331_out0;
wire  [3:0] v$_332_out1;
wire  [3:0] v$_358_out0;
wire  [3:0] v$_444_out1;
wire  [3:0] v$_454_out1;
wire  [3:0] v$_478_out0;
wire  [3:0] v$_48_out0;
wire  [3:0] v$_614_out1;
wire  [3:0] v$_727_out0;
wire  [4:0] v$4_282_out0;
wire  [4:0] v$K_13_out0;
wire  [4:0] v$_24_out1;
wire  [4:0] v$_683_out1;
wire  [5:0] v$_346_out1;
wire  [5:0] v$_633_out1;
wire  [6:0] v$NA_193_out0;
wire  [6:0] v$_354_out1;
wire  [6:0] v$_514_out0;
wire  [6:0] v$_574_out1;
wire  [7:0] v$15TO8_692_out0;
wire  [7:0] v$7TO0_476_out0;
wire  [7:0] v$C1_302_out0;
wire  [7:0] v$ZERO_34_out0;
wire  [7:0] v$_2_out0;
wire  [7:0] v$_303_out1;
wire  [7:0] v$_390_out0;
wire  [7:0] v$_390_out1;
wire  [7:0] v$_528_out0;
wire  [7:0] v$_591_out1;
wire  [7:0] v$_85_out0;
wire  [8:0] v$_338_out1;
wire  [8:0] v$_690_out1;
wire  [9:0] v$_645_out1;
wire  [9:0] v$_658_out1;
wire v$1_655_out0;
wire v$2_219_out0;
wire v$3_327_out0;
wire v$5_554_out0;
wire v$6_580_out0;
wire v$7_267_out0;
wire v$7_559_out0;
wire v$8_162_out0;
wire v$A1_135_out1;
wire v$A1_369_out1;
wire v$A1_38_out1;
wire v$ADC_153_out0;
wire v$ADC_409_out0;
wire v$ADD_451_out0;
wire v$ADD_676_out0;
wire v$AND_269_out0;
wire v$AND_5_out0;
wire v$C1_143_out0;
wire v$C1_147_out0;
wire v$C1_509_out0;
wire v$C1_585_out0;
wire v$C1_697_out0;
wire v$C2_401_out0;
wire v$C2_73_out0;
wire v$C3_539_out0;
wire v$C4_146_out0;
wire v$CIN_404_out0;
wire v$CMP_125_out0;
wire v$CMP_420_out0;
wire v$CONTEXTSAVEN_735_out0;
wire v$COUT_438_out0;
wire v$C_101_out0;
wire v$C_133_out0;
wire v$C_137_out0;
wire v$C_336_out0;
wire v$D1_500_out0;
wire v$D1_500_out1;
wire v$D1_500_out2;
wire v$D1_500_out3;
wire v$EN_166_out0;
wire v$EN_513_out0;
wire v$EN_678_out0;
wire v$EN_747_out0;
wire v$EQ1_158_out0;
wire v$EQ1_334_out0;
wire v$EQ1_483_out0;
wire v$EQ1_638_out0;
wire v$EQ1_726_out0;
wire v$EQ1_84_out0;
wire v$EQ2_326_out0;
wire v$EQ2_562_out0;
wire v$EQ2_704_out0;
wire v$EQ3_237_out0;
wire v$EQ3_556_out0;
wire v$EQ3_600_out0;
wire v$EQ4_365_out0;
wire v$EQ5_191_out0;
wire v$EQ6_479_out0;
wire v$EQ7_53_out0;
wire v$EQ8_495_out0;
wire v$EQ_105_out0;
wire v$EQ_178_out0;
wire v$EQ_292_out0;
wire v$EQ_443_out0;
wire v$EXEC1_18_out0;
wire v$EXEC1_299_out0;
wire v$EXEC1_381_out0;
wire v$EXEC1_459_out0;
wire v$EXEC1_494_out0;
wire v$EXEC1_534_out0;
wire v$EXEC1_553_out0;
wire v$EXEC2_197_out0;
wire v$EXEC2_203_out0;
wire v$EXEC2_275_out0;
wire v$EXEC2_293_out0;
wire v$EXEC2_502_out0;
wire v$EXEC2_549_out0;
wire v$EXEC2_586_out0;
wire v$EXEC2_596_out0;
wire v$EXEC2_60_out0;
wire v$EXEC2_63_out0;
wire v$EXEC2_699_out0;
wire v$FETCH_289_out0;
wire v$FETCH_364_out0;
wire v$FETCH_493_out0;
wire v$G10_281_out0;
wire v$G10_371_out0;
wire v$G10_413_out0;
wire v$G10_428_out0;
wire v$G10_708_out0;
wire v$G11_10_out0;
wire v$G11_159_out0;
wire v$G11_261_out0;
wire v$G11_575_out0;
wire v$G12_424_out0;
wire v$G12_717_out0;
wire v$G12_719_out0;
wire v$G13_246_out0;
wire v$G13_37_out0;
wire v$G14_227_out0;
wire v$G14_32_out0;
wire v$G15_291_out0;
wire v$G16_223_out0;
wire v$G1_103_out0;
wire v$G1_113_out0;
wire v$G1_130_out0;
wire v$G1_144_out0;
wire v$G1_233_out0;
wire v$G1_236_out0;
wire v$G1_497_out0;
wire v$G1_62_out0;
wire v$G2_213_out0;
wire v$G2_277_out0;
wire v$G2_373_out0;
wire v$G2_447_out0;
wire v$G2_499_out0;
wire v$G2_569_out0;
wire v$G2_689_out0;
wire v$G2_81_out0;
wire v$G3_0_out0;
wire v$G3_273_out0;
wire v$G3_295_out0;
wire v$G3_431_out0;
wire v$G3_448_out0;
wire v$G3_595_out0;
wire v$G4_286_out0;
wire v$G4_582_out0;
wire v$G4_613_out0;
wire v$G4_623_out0;
wire v$G4_646_out0;
wire v$G5_230_out0;
wire v$G5_466_out0;
wire v$G5_684_out0;
wire v$G5_734_out0;
wire v$G5_83_out0;
wire v$G6_183_out0;
wire v$G6_385_out0;
wire v$G6_50_out0;
wire v$G6_593_out0;
wire v$G6_615_out0;
wire v$G7_503_out0;
wire v$G7_541_out0;
wire v$G7_651_out0;
wire v$G7_688_out0;
wire v$G7_714_out0;
wire v$G8_134_out0;
wire v$G8_345_out0;
wire v$G8_368_out0;
wire v$G8_557_out0;
wire v$G8_663_out0;
wire v$G9_167_out0;
wire v$G9_492_out0;
wire v$G9_560_out0;
wire v$G9_627_out0;
wire v$G9_713_out0;
wire v$IJUMP_160_out0;
wire v$INTERRUPT_612_out0;
wire v$INTERRUPT_8_out0;
wire v$IR15_361_out0;
wire v$IR15_36_out0;
wire v$JEQN_262_out0;
wire v$JEQN_396_out0;
wire v$JMIN_23_out0;
wire v$JMIN_342_out0;
wire v$JMPN_122_out0;
wire v$JMPN_226_out0;
wire v$JMP_244_out0;
wire v$L_189_out0;
wire v$MI_154_out0;
wire v$MI_225_out0;
wire v$MI_421_out0;
wire v$MI_662_out0;
wire v$MOV_239_out0;
wire v$MOV_496_out0;
wire v$MUX15_632_out0;
wire v$MUX16_538_out0;
wire v$MUX17_208_out0;
wire v$MUX18_682_out0;
wire v$MUX2_188_out0;
wire v$MUX2_308_out0;
wire v$MUX2_441_out0;
wire v$MUX2_661_out0;
wire v$MUX3_455_out0;
wire v$MUX3_636_out0;
wire v$MUX3_666_out0;
wire v$MUX4_405_out0;
wire v$MUX5_296_out0;
wire v$MUX6_380_out0;
wire v$MUX7_319_out0;
wire v$MUX8_311_out0;
wire v$MUX8_379_out0;
wire v$NA_644_out0;
wire v$NOR_432_out0;
wire v$NOTUSED_674_out0;
wire v$P_102_out0;
wire v$RAMWEN_422_out0;
wire v$READREQ_374_out0;
wire v$RET_243_out0;
wire v$RET_252_out0;
wire v$RET_274_out0;
wire v$RET_278_out0;
wire v$RET_449_out0;
wire v$RET_568_out0;
wire v$RET_584_out0;
wire v$RET_74_out0;
wire v$RET_79_out0;
wire v$SBC_247_out0;
wire v$SBC_640_out0;
wire v$SEL2_149_out0;
wire v$STALL_305_out0;
wire v$STALL_536_out0;
wire v$STALL_605_out0;
wire v$STALL_611_out0;
wire v$STALL_635_out0;
wire v$STALL_695_out0;
wire v$STALL_741_out0;
wire v$STORESHADOW_195_out0;
wire v$STORESHADOW_220_out0;
wire v$STORESHADOW_301_out0;
wire v$STORESHADOW_462_out0;
wire v$STORESHADOW_471_out0;
wire v$STORESHADOW_679_out0;
wire v$STORESHADOW_77_out0;
wire v$STORESHADOW_96_out0;
wire v$STP_204_out0;
wire v$STP_313_out0;
wire v$STP_603_out0;
wire v$SUB_316_out0;
wire v$SUB_450_out0;
wire v$S_445_out0;
wire v$S_599_out0;
wire v$TST_136_out0;
wire v$TST_92_out0;
wire v$U_200_out0;
wire v$U_6_out0;
wire v$WEN3_107_out0;
wire v$WENALU_352_out0;
wire v$WENALU_739_out0;
wire v$WENLDST_121_out0;
wire v$WENLDST_39_out0;
wire v$WENRAM_703_out0;
wire v$WRITEREQ_259_out0;
wire v$W_229_out0;
wire v$X_578_out0;
wire v$_150_out0;
wire v$_151_out0;
wire v$_151_out1;
wire v$_155_out0;
wire v$_175_out0;
wire v$_175_out1;
wire v$_184_out0;
wire v$_184_out1;
wire v$_1_out0;
wire v$_202_out0;
wire v$_207_out0;
wire v$_211_out0;
wire v$_21_out0;
wire v$_231_out0;
wire v$_231_out1;
wire v$_24_out0;
wire v$_25_out0;
wire v$_270_out0;
wire v$_270_out1;
wire v$_272_out0;
wire v$_287_out1;
wire v$_303_out0;
wire v$_332_out0;
wire v$_338_out0;
wire v$_346_out0;
wire v$_350_out0;
wire v$_354_out0;
wire v$_378_out0;
wire v$_387_out0;
wire v$_411_out0;
wire v$_423_out0;
wire v$_423_out1;
wire v$_470_out1;
wire v$_501_out0;
wire v$_504_out0;
wire v$_504_out1;
wire v$_514_out1;
wire v$_552_out0;
wire v$_572_out0;
wire v$_572_out1;
wire v$_574_out0;
wire v$_57_out0;
wire v$_57_out1;
wire v$_589_out0;
wire v$_589_out1;
wire v$_591_out0;
wire v$_608_out0;
wire v$_608_out1;
wire v$_633_out0;
wire v$_645_out0;
wire v$_654_out0;
wire v$_658_out0;
wire v$_672_out0;
wire v$_683_out0;
wire v$_690_out0;
wire v$_694_out1;
wire v$_698_out0;
wire v$_709_out0;
wire v$_709_out1;
wire v$_733_out0;
wire v$_88_out0;
wire v$_99_out0;
wire v$interruptatexec2_535_out0;
wire v$interruptatexec2_668_out0;
wire v$interruptatexec2_686_out0;

always @(posedge clk) v$FF1_14_out0 <= v$STALL_305_out0;
always @(posedge clk) v$REG1_43_out0 <= v$G10_428_out0 ? v$MUX5_366_out0 : v$REG1_43_out0;
always @(posedge clk) v$REG3_65_out0 <= v$STORESHADOW_96_out0 ? v$G4_582_out0 : v$REG3_65_out0;
always @(posedge clk) v$REG2_86_out0 <= v$interruptatexec2_668_out0 ? v$MUX7_592_out0 : v$REG2_86_out0;
always @(posedge clk) v$REG1_164_out0 <= v$MUX16_538_out0 ? v$MUX12_15_out0 : v$REG1_164_out0;
always @(posedge clk) v$FF1_186_out0 <= v$_501_out0;
always @(posedge clk) v$FF1_192_out0 <= v$_589_out0;
always @(posedge clk) v$REG4_215_out0 <= v$CONTEXTSAVEN_735_out0 ? v$R3_232_out0 : v$REG4_215_out0;
always @(posedge clk) v$REG2_235_out0 <= v$STORESHADOW_96_out0 ? v$G1_233_out0 : v$REG2_235_out0;
always @(posedge clk) v$FF1_248_out0 <= v$STALL_635_out0;
always @(posedge clk) v$REG3_263_out0 <= v$CONTEXTSAVEN_735_out0 ? v$R2_391_out0 : v$REG3_263_out0;
always @(posedge clk) v$FF2_325_out0 <= v$STORESHADOW_195_out0 ? v$FF1_386_out0 : v$FF2_325_out0;
always @(posedge clk) v$REG1_339_out0 <= v$CONTEXTSAVEN_735_out0 ? v$R0_124_out0 : v$REG1_339_out0;
always @(posedge clk) v$REG2_355_out0 <= v$CONTEXTSAVEN_735_out0 ? v$R1_588_out0 : v$REG2_355_out0;
always @(posedge clk) v$REG3_383_out0 <= v$MUX18_682_out0 ? v$MUX14_198_out0 : v$REG3_383_out0;
always @(posedge clk) v$FF1_386_out0 <= v$G11_10_out0 ? v$MUX8_311_out0 : v$FF1_386_out0;
always @(posedge clk) v$REG5_394_out0 <= v$G10_413_out0 ? v$RM_392_out0 : v$REG5_394_out0;
always @(posedge clk) v$FF4_416_out0 <= v$_184_out1;
always @(posedge clk) v$REG1_434_out0 <= v$EXEC2_293_out0 ? v$ALUOUT_174_out0 : v$REG1_434_out0;
always @(posedge clk) v$FF2_437_out0 <= v$G14_227_out0 ? v$INTERRUPT_8_out0 : v$FF2_437_out0;
always @(posedge clk) v$REG1_485_out0 <= v$G2_277_out0 ? v$RAMDOUT_337_out0 : v$REG1_485_out0;
always @(posedge clk) v$FF1_564_out0 <= v$G4_646_out0 ? v$INTERRUPT_8_out0 : v$FF1_564_out0;
always @(posedge clk) v$FF2_570_out0 <= v$_589_out1;
always @(posedge clk) v$FF2_601_out0 <= v$_287_out1;
always @(posedge clk) v$FF3_606_out0 <= v$_184_out0;
always @(posedge clk) v$REG0_622_out0 <= v$MUX15_632_out0 ? v$MUX11_165_out0 : v$REG0_622_out0;
always @(posedge clk) v$REG4_660_out0 <= v$EXEC2_293_out0 ? v$ALUOUT_174_out0 : v$REG4_660_out0;
always @(posedge clk) v$REG2_665_out0 <= v$MUX17_208_out0 ? v$MUX13_548_out0 : v$REG2_665_out0;
assign v$C2_743_out0 = 16'hffff;
assign v$C1_697_out0 = 1'h0;
assign v$C1_585_out0 = 1'h0;
assign v$C1_540_out0 = 2'h0;
assign v$C3_539_out0 = 1'h0;
assign v$C1_509_out0 = 1'h1;
assign v$C1_486_out0 = 4'h0;
assign v$ROR_430_out0 = 2'h3;
assign v$C4_406_out0 = 12'h20;
assign v$C2_401_out0 = 1'h0;
assign v$C1_302_out0 = 8'h0;
assign v$C1_245_out0 = 12'h0;
assign v$C1_209_out0 = 12'h0;
assign v$C3_179_out0 = 16'h0;
assign v$C1_147_out0 = 1'h1;
assign v$C4_146_out0 = 1'h1;
assign v$C1_143_out0 = 1'h1;
assign v$C1_141_out0 = 11'h0;
assign v$C1_97_out0 = 16'h0;
assign v$C2_73_out0 = 1'h0;
assign v$C4_46_out0 = 16'hffff;
assign v$INTERRUPT_8_out0 = v$INTERRUPT_418_out0;
assign v$ZERO_34_out0 = v$C1_302_out0;
assign v$R0_106_out0 = v$REG0_622_out0;
assign v$PC1_115_out0 = v$REG1_43_out0;
assign v$R0_124_out0 = v$REG0_622_out0;
assign v$C_133_out0 = v$FF2_325_out0;
assign v$R0S_148_out0 = v$REG1_339_out0;
assign v$_196_out0 = { v$FF3_606_out0,v$FF4_416_out0 };
assign v$R3_232_out0 = v$REG3_383_out0;
assign v$G11_261_out0 = ! v$FF1_248_out0;
assign v$R2_264_out0 = v$REG2_665_out0;
assign v$PRIORITY_333_out0 = v$FF2_437_out0;
assign v$R3_363_out0 = v$REG3_383_out0;
assign v$RAMDOUT_367_out0 = v$PCORROM_461_out0;
assign {v$A1_369_out1,v$A1_369_out0 } = v$REG1_43_out0 + v$C1_209_out0 + v$C1_143_out0;
assign v$R2_391_out0 = v$REG2_665_out0;
assign v$STOREDPC_415_out0 = v$REG2_86_out0;
assign v$ZERO_426_out0 = v$C1_486_out0;
assign v$ZERO_439_out0 = v$C1_540_out0;
assign v$G3_448_out0 = ! v$FF1_14_out0;
assign v$R2S_467_out0 = v$REG3_263_out0;
assign v$_480_out0 = { v$FF1_192_out0,v$FF2_570_out0 };
assign v$R1_490_out0 = v$REG1_164_out0;
assign v$EQ2_562_out0 = v$REG1_434_out0 == 16'h0;
assign v$R1_588_out0 = v$REG1_164_out0;
assign v$PC_590_out0 = v$REG1_43_out0;
assign v$R3S_648_out0 = v$REG4_215_out0;
assign v$1_655_out0 = v$REG4_660_out0[15:15];
assign v$R1S_669_out0 = v$REG2_355_out0;
assign v$SHIFTPREVIOUS_187_out0 = v$_196_out0;
assign v$RAMDOUT_337_out0 = v$RAMDOUT_367_out0;
assign v$RAMDOUT_356_out0 = v$RAMDOUT_367_out0;
assign v$Q_517_out0 = v$_480_out0;
assign v$X_578_out0 = v$A1_369_out1;
assign v$STOREDPC_718_out0 = v$STOREDPC_415_out0;
assign v$EQ3_237_out0 = v$SHIFTPREVIOUS_187_out0 == 2'h2;
assign v$EQ2_326_out0 = v$SHIFTPREVIOUS_187_out0 == 2'h1;
assign v$EQ3_600_out0 = v$Q_517_out0 == 2'h2;
assign v$EQ1_638_out0 = v$Q_517_out0 == 2'h1;
assign v$RAMDOUT_639_out0 = v$RAMDOUT_356_out0;
assign v$EQ2_704_out0 = v$Q_517_out0 == 2'h0;
assign v$Q_729_out0 = v$Q_517_out0;
assign v$_211_out0 = v$Q_729_out0[1:1];
assign v$G1_236_out0 = v$EQ2_326_out0 && v$FF2_601_out0;
assign v$RAMDOUT_254_out0 = v$RAMDOUT_639_out0;
assign v$FETCH_364_out0 = v$EQ2_704_out0;
assign v$EXEC1_459_out0 = v$EQ1_638_out0;
assign v$_552_out0 = v$Q_729_out0[0:0];
assign v$G2_569_out0 = v$FF1_186_out0 && v$EQ3_237_out0;
assign v$EXEC2_699_out0 = v$EQ3_600_out0;
assign v$EXEC1_18_out0 = v$EXEC1_459_out0;
assign v$G1_103_out0 = ! v$_211_out0;
assign v$EXEC2_203_out0 = v$EXEC2_699_out0;
assign v$FETCH_289_out0 = v$FETCH_364_out0;
assign v$EXEC2_63_out0 = v$EXEC2_203_out0;
assign v$FETCH_493_out0 = v$FETCH_289_out0;
assign v$EXEC1_534_out0 = v$EXEC1_18_out0;
assign v$G3_295_out0 = v$EXEC2_63_out0 && v$FF1_564_out0;
assign v$EXEC1_299_out0 = v$EXEC1_534_out0;
assign v$EXEC2_502_out0 = v$EXEC2_63_out0;
assign v$EXEC2_549_out0 = v$EXEC2_63_out0;
assign v$EXEC1_553_out0 = v$EXEC1_534_out0;
assign v$G8_557_out0 = v$EXEC2_63_out0 && v$INTERRUPT_8_out0;
assign v$G6_615_out0 = v$INTERRUPT_8_out0 && v$FETCH_493_out0;
assign v$G4_646_out0 = v$INTERRUPT_8_out0 || v$FETCH_493_out0;
assign v$G2_689_out0 = v$FF1_564_out0 && v$FETCH_493_out0;
assign v$EXEC2_197_out0 = v$EXEC2_549_out0;
assign v$EXEC2_275_out0 = v$EXEC2_502_out0;
assign v$G2_277_out0 = v$EXEC1_299_out0 && v$G3_448_out0;
assign v$EXEC1_494_out0 = v$EXEC1_553_out0;
assign v$G7_688_out0 = v$G8_557_out0 || v$G3_295_out0;
assign v$G5_734_out0 = v$G2_689_out0 || v$G6_615_out0;
assign v$EXEC2_60_out0 = v$EXEC2_197_out0;
assign v$STORESHADOW_301_out0 = v$G5_734_out0;
assign v$MUX1_349_out0 = v$G2_277_out0 ? v$RAMDOUT_337_out0 : v$REG1_485_out0;
assign v$EXEC1_381_out0 = v$EXEC1_494_out0;
assign v$interruptatexec2_535_out0 = v$G7_688_out0;
assign v$EXEC2_596_out0 = v$EXEC2_197_out0;
assign v$IR_27_out0 = v$MUX1_349_out0;
assign v$STORESHADOW_77_out0 = v$STORESHADOW_301_out0;
assign v$EXEC2_293_out0 = v$EXEC2_60_out0;
assign v$G10_413_out0 = v$EXEC1_381_out0 && v$G11_261_out0;
assign v$STORESHADOW_471_out0 = v$STORESHADOW_301_out0;
assign v$EXEC2_586_out0 = v$EXEC2_596_out0;
assign v$INTERRUPT_612_out0 = v$interruptatexec2_535_out0;
assign v$_614_out0 = v$MUX1_349_out0[11:0];
assign v$_614_out1 = v$MUX1_349_out0[15:4];
assign v$interruptatexec2_686_out0 = v$interruptatexec2_535_out0;
assign v$EQ7_53_out0 = v$_614_out1 == 4'h6;
assign v$STORESHADOW_96_out0 = v$STORESHADOW_471_out0;
assign v$EQ5_191_out0 = v$_614_out1 == 4'h4;
assign v$STORESHADOW_195_out0 = v$STORESHADOW_471_out0;
assign v$STORESHADOW_220_out0 = v$STORESHADOW_471_out0;
assign v$STORESHADOW_462_out0 = v$STORESHADOW_77_out0;
assign v$EQ6_479_out0 = v$_614_out1 == 4'h5;
assign v$EQ8_495_out0 = v$_614_out1 == 4'h7;
assign v$interruptatexec2_668_out0 = v$interruptatexec2_686_out0;
assign v$IR110_675_out0 = v$_614_out0;
assign v$IR16_716_out0 = v$IR_27_out0;
assign v$EQ1_726_out0 = v$_614_out1 == 4'h3;
assign v$SEL1_64_out0 = v$IR16_716_out0[15:12];
assign v$G1_144_out0 = v$INTERRUPT_612_out0 || v$EQ5_191_out0;
assign v$SEL2_149_out0 = v$IR16_716_out0[9:9];
assign v$JEQN_262_out0 = v$EQ7_53_out0;
assign v$G3_273_out0 = v$STORESHADOW_462_out0 || v$interruptatexec2_668_out0;
assign v$STP_313_out0 = v$EQ8_495_out0;
assign v$JMIN_342_out0 = v$EQ6_479_out0;
assign v$IR12_436_out0 = v$IR110_675_out0;
assign v$IR_526_out0 = v$IR16_716_out0;
assign v$RET_568_out0 = v$EQ1_726_out0;
assign v$STORESHADOW_679_out0 = v$STORESHADOW_220_out0;
assign v$3_4_out0 = v$IR_526_out0[1:0];
assign v$8_11_out0 = v$IR_526_out0[11:10];
assign v$JMIN_23_out0 = v$JMIN_342_out0;
assign v$IJUMP_160_out0 = v$G3_273_out0;
assign v$JMPN_226_out0 = v$G1_144_out0;
assign v$IR_297_out0 = v$IR_526_out0;
assign v$EQ1_334_out0 = v$SEL1_64_out0 == 4'h0;
assign v$JEQN_396_out0 = v$JEQN_262_out0;
assign v$7_559_out0 = v$IR_526_out0[15:15];
assign v$G9_560_out0 = v$SEL2_149_out0 && v$EXEC1_534_out0;
assign v$RET_584_out0 = v$RET_568_out0;
assign v$1_597_out0 = v$IR_526_out0[14:12];
assign v$STP_603_out0 = v$STP_313_out0;
assign v$N_681_out0 = v$IR12_436_out0;
assign v$CONTEXTSAVEN_735_out0 = v$STORESHADOW_679_out0;
assign v$IR15_36_out0 = v$7_559_out0;
assign v$5_71_out0 = v$IR_297_out0[7:4];
assign v$RET_74_out0 = v$RET_584_out0;
assign v$OP_110_out0 = v$1_597_out0;
assign v$JMPN_122_out0 = v$JMPN_226_out0;
assign v$9_131_out0 = v$IR_297_out0[3:2];
assign v$M_138_out0 = v$3_4_out0;
assign v$STP_204_out0 = v$STP_603_out0;
assign v$2_219_out0 = v$IR_297_out0[8:8];
assign v$G14_227_out0 = v$INTERRUPT_8_out0 || v$RET_584_out0;
assign v$RET_243_out0 = v$RET_584_out0;
assign v$4_282_out0 = v$IR_297_out0[4:0];
assign v$IR_330_out0 = v$IR_297_out0;
assign v$D_359_out0 = v$8_11_out0;
assign v$MUX6_456_out0 = v$interruptatexec2_668_out0 ? v$C4_406_out0 : v$N_681_out0;
assign v$6_580_out0 = v$IR_297_out0[9:9];
assign v$G10_708_out0 = v$EQ1_334_out0 && v$G9_560_out0;
assign v$K_13_out0 = v$4_282_out0;
assign v$OP_58_out0 = v$OP_110_out0;
assign v$RET_79_out0 = v$RET_74_out0;
assign v$IR_94_out0 = v$IR_330_out0;
assign v$C_101_out0 = v$6_580_out0;
assign v$MUX2_112_out0 = v$EXEC2_197_out0 ? v$D_359_out0 : v$M_138_out0;
assign v$JMP_244_out0 = v$JMPN_122_out0;
assign v$SHIFT_271_out0 = v$9_131_out0;
assign v$RET_274_out0 = v$RET_243_out0;
assign v$RET_278_out0 = v$RET_74_out0;
assign v$IR15_361_out0 = v$IR15_36_out0;
assign v$READREQ_374_out0 = v$G10_708_out0;
assign v$RET_449_out0 = v$RET_74_out0;
assign v$B_464_out0 = v$5_71_out0;
assign v$AD2_581_out0 = v$M_138_out0;
assign v$S_599_out0 = v$2_219_out0;
assign v$AD1_742_out0 = v$D_359_out0;
assign v$AND_5_out0 = v$OP_58_out0 == 3'h6;
assign v$G1_62_out0 = v$EXEC2_586_out0 && v$IR15_361_out0;
assign v$B_66_out0 = v$B_464_out0;
assign v$TST_92_out0 = v$OP_58_out0 == 3'h7;
assign v$_108_out0 = { v$K_13_out0,v$C1_141_out0 };
assign v$G1_113_out0 = v$JMP_244_out0 || v$RET_243_out0;
assign v$6_116_out0 = v$IR_94_out0[1:0];
assign v$C_137_out0 = v$C_101_out0;
assign v$8_162_out0 = v$IR_94_out0[8:8];
assign v$_231_out0 = v$AD2_581_out0[0:0];
assign v$_231_out1 = v$AD2_581_out0[1:1];
assign v$RET_252_out0 = v$RET_79_out0;
assign v$7_267_out0 = v$IR_94_out0[6:6];
assign v$4_288_out0 = v$IR_94_out0[15:12];
assign v$3_327_out0 = v$IR_94_out0[7:7];
assign v$9_400_out0 = v$IR_94_out0[5:2];
assign v$ADC_409_out0 = v$OP_58_out0 == 3'h2;
assign v$CMP_420_out0 = v$OP_58_out0 == 3'h5;
assign v$_423_out0 = v$AD1_742_out0[0:0];
assign v$_423_out1 = v$AD1_742_out0[1:1];
assign v$S_445_out0 = v$S_599_out0;
assign v$SUB_450_out0 = v$OP_58_out0 == 3'h1;
assign v$ADD_451_out0 = v$OP_58_out0 == 3'h0;
assign v$2_468_out0 = v$IR_94_out0[11:10];
assign v$MOV_496_out0 = v$OP_58_out0 == 3'h4;
assign v$AD3_550_out0 = v$MUX2_112_out0;
assign v$5_554_out0 = v$IR_94_out0[9:9];
assign v$G11_575_out0 = ((v$READVALID_17_out0 && !v$READREQ_374_out0) || (!v$READVALID_17_out0) && v$READREQ_374_out0);
assign v$SBC_640_out0 = v$OP_58_out0 == 3'h3;
assign v$SR_659_out0 = v$SHIFT_271_out0;
assign v$U_6_out0 = v$7_267_out0;
assign v$G11_10_out0 = v$S_445_out0 && v$EXEC2_586_out0;
assign v$MUX4_51_out0 = v$_231_out0 ? v$R1_490_out0 : v$R0_106_out0;
assign v$D_59_out0 = v$2_468_out0;
assign v$P_102_out0 = v$3_327_out0;
assign v$B_114_out0 = v$B_66_out0;
assign v$CMP_125_out0 = v$CMP_420_out0;
assign v$TST_136_out0 = v$TST_92_out0;
assign v$ADC_153_out0 = v$ADC_409_out0;
assign v$L_189_out0 = v$5_554_out0;
assign v$MUX8_206_out0 = v$RET_252_out0 ? v$R1S_669_out0 : v$R1_490_out0;
assign v$G2_213_out0 = v$G1_113_out0 || v$G3_273_out0;
assign v$W_229_out0 = v$8_162_out0;
assign v$MOV_239_out0 = v$MOV_496_out0;
assign v$SBC_247_out0 = v$SBC_640_out0;
assign v$MUX10_266_out0 = v$RET_252_out0 ? v$R3S_648_out0 : v$R3_363_out0;
assign v$AND_269_out0 = v$AND_5_out0;
assign v$O_312_out0 = v$4_288_out0;
assign v$SUB_316_out0 = v$SUB_450_out0;
assign v$C_336_out0 = v$C_137_out0;
assign v$N_343_out0 = v$9_400_out0;
assign v$MUX7_389_out0 = v$RET_252_out0 ? v$R0S_148_out0 : v$R0_106_out0;
assign v$MUX5_498_out0 = v$_231_out0 ? v$R3_363_out0 : v$R2_264_out0;
assign v$MUX9_508_out0 = v$RET_252_out0 ? v$R2S_467_out0 : v$R2_264_out0;
assign v$M_629_out0 = v$6_116_out0;
assign v$ADD_676_out0 = v$ADD_451_out0;
assign v$_733_out0 = v$B_66_out0[0:0];
assign v$_733_out1 = v$B_66_out0[3:3];
assign v$MUX1_3_out0 = v$C_336_out0 ? v$ROR_430_out0 : v$SR_659_out0;
assign v$R1S_29_out0 = v$MUX8_206_out0;
assign v$G6_50_out0 = v$EXEC1_381_out0 && v$W_229_out0;
assign v$EQ1_84_out0 = v$O_312_out0 == 4'h6;
assign v$G8_134_out0 = v$SUB_316_out0 || v$CMP_125_out0;
assign v$R0S_140_out0 = v$MUX7_389_out0;
assign v$R2S_161_out0 = v$MUX9_508_out0;
assign v$MUX6_170_out0 = v$_231_out1 ? v$MUX5_498_out0 : v$MUX4_51_out0;
assign v$MUX2_188_out0 = v$ADD_676_out0 ? v$C2_401_out0 : v$FF1_386_out0;
assign v$U_200_out0 = v$U_6_out0;
assign v$G5_230_out0 = ! v$MOV_239_out0;
assign v$B_241_out0 = v$B_114_out0;
assign v$R3TEST_242_out0 = v$MUX10_266_out0;
assign v$_350_out0 = v$_733_out1[0:0];
assign v$_350_out1 = v$_733_out1[2:2];
assign v$EQ4_365_out0 = v$O_312_out0 == 4'h0;
assign v$G2_373_out0 = ! v$C_336_out0;
assign v$G3_431_out0 = v$EXEC2_293_out0 && v$L_189_out0;
assign v$G2_447_out0 = ! v$L_189_out0;
assign v$EQ1_483_out0 = v$B_114_out0 == 4'h0;
assign v$G9_492_out0 = !(v$CMP_125_out0 || v$TST_136_out0);
assign v$G2_499_out0 = v$SUB_316_out0 || v$SBC_247_out0;
assign v$EQ3_556_out0 = v$O_312_out0 == 4'h5;
assign v$G3_595_out0 = v$ADD_676_out0 || v$ADC_153_out0;
assign v$R3S_650_out0 = v$MUX10_266_out0;
assign v$G8_663_out0 = v$L_189_out0 && v$EXEC2_293_out0;
assign v$N_715_out0 = v$N_343_out0;
assign v$G12_719_out0 = v$AND_269_out0 || v$TST_136_out0;
assign v$DOUT2_117_out0 = v$MUX6_170_out0;
assign v$EQ1_158_out0 = v$B_241_out0 == 4'h0;
assign v$EN_166_out0 = v$_350_out0;
assign v$MUX1_194_out0 = v$_423_out0 ? v$R1S_29_out0 : v$R0S_140_out0;
assign v$G1_233_out0 = v$EQ1_84_out0 && v$EQ2_562_out0;
assign v$R0TEST_283_out0 = v$R0S_140_out0;
assign v$_320_out0 = { v$N_715_out0,v$C1_245_out0 };
assign v$MUX2_360_out0 = v$_423_out0 ? v$R3S_650_out0 : v$R2S_161_out0;
assign v$SR_414_out0 = v$MUX1_3_out0;
assign v$NOR_432_out0 = v$G9_492_out0;
assign v$MUX2_441_out0 = v$U_200_out0 ? v$C3_539_out0 : v$C4_146_out0;
assign v$G5_466_out0 = v$G6_50_out0 || v$G3_431_out0;
assign v$G1_497_out0 = v$G2_373_out0 && v$_733_out0;
assign v$R1TEST_551_out0 = v$R1S_29_out0;
assign v$_572_out0 = v$_350_out1[0:0];
assign v$_572_out1 = v$_350_out1[1:1];
assign v$G4_582_out0 = v$1_655_out0 && v$EQ3_556_out0;
assign v$R2TEST_583_out0 = v$R2S_161_out0;
assign v$MUX3_636_out0 = v$G8_134_out0 ? v$C1_509_out0 : v$MUX2_188_out0;
assign v$G7_651_out0 = v$G2_499_out0 || v$CMP_125_out0;
assign v$G9_713_out0 = v$EXEC2_293_out0 && v$G2_447_out0;
assign v$R3TEST_732_out0 = v$R3TEST_242_out0;
assign v$WENLDST_39_out0 = v$G5_466_out0;
assign v$MUX3_42_out0 = v$_423_out1 ? v$MUX2_360_out0 : v$MUX1_194_out0;
assign v$SR_104_out0 = v$SR_414_out0;
assign v$R2TEST_152_out0 = v$R2TEST_583_out0;
assign v$SHIFT_182_out0 = v$SR_414_out0;
assign v$XOR1_253_out0 = v$_320_out0 ^ v$C2_743_out0;
assign v$G10_281_out0 = v$G1_62_out0 && v$NOR_432_out0;
assign v$SR_317_out0 = v$SR_414_out0;
assign v$R1TEST_376_out0 = v$R1TEST_551_out0;
assign v$CIN_404_out0 = v$MUX3_636_out0;
assign v$MUX4_405_out0 = v$RET_449_out0 ? v$REG2_235_out0 : v$G1_233_out0;
assign v$EN_513_out0 = v$G1_497_out0;
assign v$SR_537_out0 = v$SR_414_out0;
assign v$MUX1_547_out0 = v$G7_651_out0 ? v$C4_46_out0 : v$C3_179_out0;
assign v$SR_565_out0 = v$SR_414_out0;
assign v$G4_613_out0 = v$G7_651_out0 || v$G3_595_out0;
assign v$RM_620_out0 = v$DOUT2_117_out0;
assign v$MUX2_661_out0 = v$RET_449_out0 ? v$REG3_65_out0 : v$G4_582_out0;
assign v$EN_678_out0 = v$_572_out0;
assign v$RM_685_out0 = v$DOUT2_117_out0;
assign v$R3_693_out0 = v$R3TEST_732_out0;
assign v$R0TEST_700_out0 = v$R0TEST_283_out0;
assign v$G7_714_out0 = v$EQ4_365_out0 && v$G9_713_out0;
assign v$EN_747_out0 = v$_572_out1;
assign v$_57_out0 = v$SR_565_out0[0:0];
assign v$_57_out1 = v$SR_565_out0[1:1];
assign v$DOUT1_98_out0 = v$MUX3_42_out0;
assign v$EQ_105_out0 = v$MUX4_405_out0;
assign v$WENLDST_121_out0 = v$WENLDST_39_out0;
assign v$_151_out0 = v$SR_104_out0[0:0];
assign v$_151_out1 = v$SR_104_out0[1:1];
assign v$_184_out0 = v$SHIFT_182_out0[0:0];
assign v$_184_out1 = v$SHIFT_182_out0[1:1];
assign v$RM_210_out0 = v$RM_685_out0;
assign v$_270_out0 = v$SR_317_out0[0:0];
assign v$_270_out1 = v$SR_317_out0[1:1];
assign v$R3_276_out0 = v$R3_693_out0;
assign v$G6_385_out0 = v$G4_613_out0 && v$G5_230_out0;
assign v$RM_392_out0 = v$RM_685_out0;
assign v$MUX1_393_out0 = v$U_200_out0 ? v$_320_out0 : v$XOR1_253_out0;
assign v$MI_421_out0 = v$MUX2_661_out0;
assign v$RAMWEN_422_out0 = v$G7_714_out0;
assign v$MUX1_489_out0 = v$C_137_out0 ? v$_108_out0 : v$RM_620_out0;
assign v$_504_out0 = v$SR_537_out0[0:0];
assign v$_504_out1 = v$SR_537_out0[1:1];
assign v$R2_529_out0 = v$R2TEST_152_out0;
assign v$R1_561_out0 = v$R1TEST_376_out0;
assign v$R0_571_out0 = v$R0TEST_700_out0;
assign v$WENALU_739_out0 = v$G10_281_out0;
assign v$EQ_178_out0 = v$EQ_105_out0;
assign v$R3_251_out0 = v$R3_276_out0;
assign v$RD_260_out0 = v$DOUT1_98_out0;
assign v$RM_284_out0 = v$RM_210_out0;
assign v$SHIFTIN_300_out0 = v$MUX1_489_out0;
assign v$WENALU_352_out0 = v$WENALU_739_out0;
assign v$R1_375_out0 = v$R1_561_out0;
assign v$MUX5_403_out0 = v$G10_413_out0 ? v$RM_392_out0 : v$REG5_394_out0;
assign v$R0_519_out0 = v$R0_571_out0;
assign v$MI_662_out0 = v$MI_421_out0;
assign v$R2_687_out0 = v$R2_529_out0;
assign v$WENRAM_703_out0 = v$RAMWEN_422_out0;
assign v$RM_142_out0 = v$MUX5_403_out0;
assign v$MI_154_out0 = v$MI_662_out0;
assign v$RDOUT_216_out0 = v$RD_260_out0;
assign v$IN_222_out0 = v$SHIFTIN_300_out0;
assign v$WRITEREQ_259_out0 = v$WENRAM_703_out0;
assign v$EQ_292_out0 = v$EQ_178_out0;
assign v$R2_370_out0 = v$R2_687_out0;
assign v$R0_525_out0 = v$R0_519_out0;
assign v$OP1_555_out0 = v$RD_260_out0;
assign v$MUX3_666_out0 = v$IR15_36_out0 ? v$WENALU_352_out0 : v$WENLDST_121_out0;
assign v$IN_667_out0 = v$SHIFTIN_300_out0;
assign v$R1_691_out0 = v$R1_375_out0;
assign v$RDOUT_33_out0 = v$RDOUT_216_out0;
assign v$WEN3_107_out0 = v$MUX3_666_out0;
assign v$OP1_176_out0 = v$OP1_555_out0;
assign v$MI_225_out0 = v$MI_154_out0;
assign v$IN_384_out0 = v$IN_667_out0;
assign v$MUX3_427_out0 = v$EQ1_483_out0 ? v$IN_222_out0 : v$C1_97_out0;
assign v$EQ_443_out0 = v$EQ_292_out0;
assign v$RM_458_out0 = v$RM_142_out0;
assign v$G12_717_out0 = ((v$WRITEREQ_259_out0 && !v$WRITECOMPLETE_55_out0) || (!v$WRITEREQ_259_out0) && v$WRITECOMPLETE_55_out0);
assign v$G13_37_out0 = v$G11_575_out0 || v$G12_717_out0;
assign v$_99_out0 = v$IN_384_out0[0:0];
assign v$_99_out1 = v$IN_384_out0[15:15];
assign {v$A1_135_out1,v$A1_135_out0 } = v$RM_458_out0 + v$MUX1_393_out0 + v$MUX2_441_out0;
assign v$G6_183_out0 = v$EQ_443_out0 || v$MI_225_out0;
assign v$G4_286_out0 = v$EQ_443_out0 || v$IJUMP_160_out0;
assign v$IN_307_out0 = v$MUX3_427_out0;
assign v$_470_out0 = v$IN_384_out0[14:0];
assign v$_470_out1 = v$IN_384_out0[15:1];
assign v$D1_500_out0 = (v$AD3_550_out0 == 2'b00) ? v$WEN3_107_out0 : 1'h0;
assign v$D1_500_out1 = (v$AD3_550_out0 == 2'b01) ? v$WEN3_107_out0 : 1'h0;
assign v$D1_500_out2 = (v$AD3_550_out0 == 2'b10) ? v$WEN3_107_out0 : 1'h0;
assign v$D1_500_out3 = (v$AD3_550_out0 == 2'b11) ? v$WEN3_107_out0 : 1'h0;
assign v$A_656_out0 = v$OP1_176_out0;
assign v$G5_684_out0 = v$MI_225_out0 || v$IJUMP_160_out0;
assign v$_20_out0 = { v$_99_out1,v$_99_out0 };
assign v$MUX17_208_out0 = v$RET_252_out0 ? v$C1_147_out0 : v$D1_500_out2;
assign v$_224_out0 = { v$_99_out1,v$_470_out1 };
assign v$IN_310_out0 = v$IN_307_out0;
assign v$G8_345_out0 = v$G4_286_out0 || v$G5_684_out0;
assign v$_395_out0 = { v$_99_out1,v$C2_73_out0 };
assign v$RMN_452_out0 = v$A1_135_out0;
assign v$_510_out0 = { v$C1_697_out0,v$_470_out0 };
assign v$MUX16_538_out0 = v$RET_252_out0 ? v$C1_147_out0 : v$D1_500_out1;
assign v$MUX7_592_out0 = v$G6_183_out0 ? v$N_681_out0 : v$A1_369_out0;
assign v$MUX15_632_out0 = v$RET_252_out0 ? v$C1_147_out0 : v$D1_500_out0;
assign v$_672_out0 = v$A_656_out0[0:0];
assign v$_672_out1 = v$A_656_out0[15:15];
assign v$NOTUSED_674_out0 = v$A1_135_out1;
assign v$MUX18_682_out0 = v$RET_252_out0 ? v$C1_147_out0 : v$D1_500_out3;
assign v$STALL_741_out0 = v$G13_37_out0;
assign v$ASR_76_out0 = v$_224_out0;
assign v$RMN_95_out0 = v$RMN_452_out0;
assign v$ROR_201_out0 = v$_20_out0;
assign v$_207_out0 = v$_672_out1[0:0];
assign v$_207_out1 = v$_672_out1[14:14];
assign v$_287_out0 = v$IN_310_out0[14:0];
assign v$_287_out1 = v$IN_310_out0[15:1];
assign v$STALL_305_out0 = v$STALL_741_out0;
assign v$_501_out0 = v$IN_310_out0[0:0];
assign v$_501_out1 = v$IN_310_out0[15:15];
assign v$LSL_515_out0 = v$_510_out0;
assign v$STALL_536_out0 = v$STALL_741_out0;
assign v$G7_541_out0 = v$G2_213_out0 || v$G8_345_out0;
assign v$STALL_605_out0 = v$STALL_741_out0;
assign v$STALL_611_out0 = v$STALL_741_out0;
assign v$LSR_677_out0 = v$_395_out0;
assign v$MUX3_54_out0 = v$_504_out1 ? v$ROR_201_out0 : v$LSR_677_out0;
assign v$_69_out0 = { v$G1_236_out0,v$_287_out0 };
assign v$MUX2_87_out0 = v$G7_541_out0 ? v$MUX6_456_out0 : v$A1_369_out0;
assign v$_150_out0 = v$_207_out1[0:0];
assign v$_150_out1 = v$_207_out1[13:13];
assign v$MUX2_256_out0 = v$_504_out1 ? v$ASR_76_out0 : v$LSL_515_out0;
assign v$MUX3_442_out0 = v$G8_663_out0 ? v$RAMDOUT_254_out0 : v$RMN_95_out0;
assign v$MUX1_512_out0 = v$P_102_out0 ? v$RMN_95_out0 : v$RM_142_out0;
assign v$G9_627_out0 = ! v$STALL_605_out0;
assign v$STALL_635_out0 = v$STALL_611_out0;
assign v$STALL_695_out0 = v$STALL_536_out0;
assign v$_728_out0 = { v$_501_out1,v$G2_569_out0 };
assign v$MUX4_49_out0 = v$_504_out0 ? v$MUX3_54_out0 : v$MUX2_256_out0;
assign v$MSL_68_out0 = v$_69_out0;
assign v$MUX4_89_out0 = v$STP_204_out0 ? v$PC_590_out0 : v$MUX2_87_out0;
assign v$MUX5_296_out0 = v$STALL_695_out0 ? v$G1_103_out0 : v$C1_585_out0;
assign v$MUX2_308_out0 = v$STALL_695_out0 ? v$C1_585_out0 : v$G1_103_out0;
assign v$MUX7_319_out0 = v$STALL_695_out0 ? v$_211_out0 : v$C1_585_out0;
assign v$MSR_321_out0 = v$_728_out0;
assign v$EA_341_out0 = v$MUX1_512_out0;
assign v$MUX8_379_out0 = v$STALL_695_out0 ? v$C1_585_out0 : v$G1_103_out0;
assign v$_411_out0 = v$_150_out1[0:0];
assign v$_411_out1 = v$_150_out1[12:12];
assign v$G10_428_out0 = v$EXEC2_502_out0 && v$G9_627_out0;
assign v$_444_out0 = v$MUX1_512_out0[11:0];
assign v$_444_out1 = v$MUX1_512_out0[15:4];
assign v$REGDIN_446_out0 = v$MUX3_442_out0;
assign v$MUX4_28_out0 = v$_184_out0 ? v$IN_310_out0 : v$MSR_321_out0;
assign v$MUX1_168_out0 = v$EN_513_out0 ? v$MUX4_49_out0 : v$IN_384_out0;
assign v$RAMADDRMUX_173_out0 = v$_444_out0;
assign v$REGDIN_238_out0 = v$REGDIN_446_out0;
assign v$MUX5_366_out0 = v$RET_274_out0 ? v$REG2_86_out0 : v$MUX4_89_out0;
assign v$MUX6_380_out0 = v$_552_out0 ? v$MUX5_296_out0 : v$MUX8_379_out0;
assign v$MUX3_455_out0 = v$_552_out0 ? v$MUX2_308_out0 : v$MUX7_319_out0;
assign v$NOTUSED_649_out0 = v$_444_out1;
assign v$_698_out0 = v$_411_out1[0:0];
assign v$_698_out1 = v$_411_out1[11:11];
assign v$MUX3_724_out0 = v$_184_out0 ? v$MSL_68_out0 : v$IN_310_out0;
assign v$OUT_212_out0 = v$MUX1_168_out0;
assign v$MUX2_511_out0 = v$_184_out1 ? v$MUX4_28_out0 : v$MUX3_724_out0;
assign v$_577_out0 = { v$MUX6_380_out0,v$MUX3_455_out0 };
assign v$_645_out0 = v$_698_out1[0:0];
assign v$_645_out1 = v$_698_out1[10:10];
assign v$RAMADDRMUX_723_out0 = v$RAMADDRMUX_173_out0;
assign v$RAMADDRMUX_72_out0 = v$RAMADDRMUX_723_out0;
assign v$IN_412_out0 = v$OUT_212_out0;
assign v$MUX1_524_out0 = v$EQ1_158_out0 ? v$MUX2_511_out0 : v$IN_310_out0;
assign v$Q1_618_out0 = v$_577_out0;
assign v$_690_out0 = v$_645_out1[0:0];
assign v$_690_out1 = v$_645_out1[9:9];
assign v$_303_out0 = v$_690_out1[0:0];
assign v$_303_out1 = v$_690_out1[8:8];
assign v$OUT_399_out0 = v$MUX1_524_out0;
assign v$RAMADDRMUX_505_out0 = v$RAMADDRMUX_72_out0;
assign v$IN_619_out0 = v$IN_412_out0;
assign v$D_707_out0 = v$Q1_618_out0;
assign v$_129_out0 = v$IN_619_out0[13:0];
assign v$_129_out1 = v$IN_619_out0[15:2];
assign v$MUX1_531_out0 = v$FETCH_493_out0 ? v$PC1_115_out0 : v$RAMADDRMUX_505_out0;
assign v$_574_out0 = v$_303_out1[0:0];
assign v$_574_out1 = v$_303_out1[7:7];
assign v$_589_out0 = v$D_707_out0[0:0];
assign v$_589_out1 = v$D_707_out0[1:1];
assign v$_602_out0 = v$IN_619_out0[1:0];
assign v$_602_out1 = v$IN_619_out0[15:14];
assign v$_30_out0 = { v$_602_out1,v$ZERO_439_out0 };
assign v$_56_out0 = { v$_602_out1,v$_602_out0 };
assign v$_180_out0 = { v$ZERO_439_out0,v$_129_out0 };
assign v$_346_out0 = v$_574_out1[0:0];
assign v$_346_out1 = v$_574_out1[6:6];
assign v$_608_out0 = v$_129_out1[0:0];
assign v$_608_out1 = v$_129_out1[1:1];
assign v$PROGRAMADDRESS_616_out0 = v$MUX1_531_out0;
assign v$ROR_118_out0 = v$_56_out0;
assign v$_322_out0 = { v$_608_out1,v$_608_out1 };
assign v$LSR_402_out0 = v$_30_out0;
assign v$NA_644_out0 = v$_608_out0;
assign v$_683_out0 = v$_346_out1[0:0];
assign v$_683_out1 = v$_346_out1[5:5];
assign v$LSL_738_out0 = v$_180_out0;
assign v$_155_out0 = v$_683_out1[0:0];
assign v$_155_out1 = v$_683_out1[4:4];
assign v$_453_out0 = { v$_602_out1,v$_322_out0 };
assign v$MUX3_671_out0 = v$_57_out1 ? v$ROR_118_out0 : v$LSR_402_out0;
assign v$ASR_377_out0 = v$_453_out0;
assign v$_654_out0 = v$_155_out1[0:0];
assign v$_654_out1 = v$_155_out1[3:3];
assign v$_21_out0 = v$_654_out1[0:0];
assign v$_21_out1 = v$_654_out1[2:2];
assign v$MUX2_280_out0 = v$_57_out1 ? v$ASR_377_out0 : v$LSL_738_out0;
assign v$_175_out0 = v$_21_out1[0:0];
assign v$_175_out1 = v$_21_out1[1:1];
assign v$MUX4_234_out0 = v$_57_out0 ? v$MUX3_671_out0 : v$MUX2_280_out0;
assign v$MUX1_664_out0 = v$EN_166_out0 ? v$MUX4_234_out0 : v$IN_619_out0;
assign v$OUT_128_out0 = v$MUX1_664_out0;
assign v$IN_673_out0 = v$OUT_128_out0;
assign v$IN_41_out0 = v$IN_673_out0;
assign v$_358_out0 = v$IN_41_out0[3:0];
assign v$_358_out1 = v$IN_41_out0[15:12];
assign v$_454_out0 = v$IN_41_out0[11:0];
assign v$_454_out1 = v$IN_41_out0[15:4];
assign v$_78_out0 = { v$ZERO_426_out0,v$_454_out0 };
assign v$_566_out0 = { v$_358_out1,v$_358_out0 };
assign v$_567_out0 = { v$_358_out1,v$ZERO_426_out0 };
assign v$_694_out0 = v$_454_out1[2:0];
assign v$_694_out1 = v$_454_out1[3:1];
assign v$LSL_250_out0 = v$_78_out0;
assign v$_318_out0 = { v$_694_out1,v$_694_out1 };
assign v$ROR_324_out0 = v$_566_out0;
assign v$LSR_335_out0 = v$_567_out0;
assign v$NA_474_out0 = v$_694_out0;
assign v$_177_out0 = { v$_318_out0,v$_318_out0 };
assign v$MUX3_306_out0 = v$_151_out1 ? v$ROR_324_out0 : v$LSR_335_out0;
assign v$_109_out0 = { v$_358_out1,v$_177_out0 };
assign v$ASR_22_out0 = v$_109_out0;
assign v$MUX2_642_out0 = v$_151_out1 ? v$ASR_22_out0 : v$LSL_250_out0;
assign v$MUX4_127_out0 = v$_151_out0 ? v$MUX3_306_out0 : v$MUX2_642_out0;
assign v$MUX1_731_out0 = v$EN_678_out0 ? v$MUX4_127_out0 : v$IN_41_out0;
assign v$OUT_730_out0 = v$MUX1_731_out0;
assign v$IN_626_out0 = v$OUT_730_out0;
assign v$IN_120_out0 = v$IN_626_out0;
assign v$_390_out0 = v$IN_120_out0[7:0];
assign v$_390_out1 = v$IN_120_out0[15:8];
assign v$7TO0_476_out0 = v$_390_out0;
assign v$15TO8_692_out0 = v$_390_out1;
assign v$_44_out0 = { v$ZERO_34_out0,v$7TO0_476_out0 };
assign v$_457_out0 = { v$15TO8_692_out0,v$ZERO_34_out0 };
assign v$_481_out0 = { v$15TO8_692_out0,v$7TO0_476_out0 };
assign v$_514_out0 = v$15TO8_692_out0[6:0];
assign v$_514_out1 = v$15TO8_692_out0[7:1];
assign v$_123_out0 = { v$_514_out1,v$_514_out1 };
assign v$LSL_163_out0 = v$_44_out0;
assign v$NA_193_out0 = v$_514_out0;
assign v$LSR_268_out0 = v$_457_out0;
assign v$ROR_353_out0 = v$_481_out0;
assign v$_294_out0 = { v$_123_out0,v$_123_out0 };
assign v$MUX3_425_out0 = v$_270_out1 ? v$ROR_353_out0 : v$LSR_268_out0;
assign v$_2_out0 = { v$_294_out0,v$_294_out0 };
assign v$_398_out0 = { v$15TO8_692_out0,v$_2_out0 };
assign v$ASR_93_out0 = v$_398_out0;
assign v$MUX2_90_out0 = v$_270_out1 ? v$ASR_93_out0 : v$LSL_163_out0;
assign v$MUX4_156_out0 = v$_270_out0 ? v$MUX3_425_out0 : v$MUX2_90_out0;
assign v$MUX1_598_out0 = v$EN_747_out0 ? v$MUX4_156_out0 : v$IN_120_out0;
assign v$OUT_624_out0 = v$MUX1_598_out0;
assign v$MUX2_265_out0 = v$EQ1_483_out0 ? v$OUT_399_out0 : v$OUT_624_out0;
assign v$SHIFTOUT_221_out0 = v$MUX2_265_out0;
assign v$OP2_348_out0 = v$SHIFTOUT_221_out0;
assign v$OP2_388_out0 = v$OP2_348_out0;
assign v$OP2_546_out0 = v$OP2_388_out0;
assign v$OP2_257_out0 = v$OP2_546_out0;
assign v$XOR1_169_out0 = v$OP2_257_out0 ^ v$MUX1_547_out0;
assign v$B_558_out0 = v$OP2_257_out0;
assign v$_25_out0 = v$B_558_out0[0:0];
assign v$_25_out1 = v$B_558_out0[15:15];
assign {v$A1_38_out1,v$A1_38_out0 } = v$OP1_176_out0 + v$XOR1_169_out0 + v$CIN_404_out0;
assign v$_1_out0 = v$_25_out1[0:0];
assign v$_1_out1 = v$_25_out1[14:14];
assign v$G1_130_out0 = v$_672_out0 && v$_25_out0;
assign v$COUT_438_out0 = v$A1_38_out1;
assign v$1TO4_487_out0 = v$A1_38_out0;
assign v$G2_81_out0 = v$_207_out0 && v$_1_out0;
assign v$_272_out0 = v$_1_out1[0:0];
assign v$_272_out1 = v$_1_out1[13:13];
assign v$MUX8_311_out0 = v$RET_278_out0 ? v$C_133_out0 : v$COUT_438_out0;
assign v$MUX4_725_out0 = v$G6_385_out0 ? v$1TO4_487_out0 : v$OP2_257_out0;
assign v$G3_0_out0 = v$_150_out0 && v$_272_out0;
assign v$_202_out0 = v$_272_out1[0:0];
assign v$_202_out1 = v$_272_out1[12:12];
assign v$_746_out0 = { v$G1_130_out0,v$G2_81_out0 };
assign v$_387_out0 = v$_202_out1[0:0];
assign v$_387_out1 = v$_202_out1[11:11];
assign v$G4_623_out0 = v$_411_out0 && v$_202_out0;
assign v$G5_83_out0 = v$_698_out0 && v$_387_out0;
assign v$_520_out0 = { v$G3_0_out0,v$G4_623_out0 };
assign v$_658_out0 = v$_387_out1[0:0];
assign v$_658_out1 = v$_387_out1[10:10];
assign v$_331_out0 = { v$_746_out0,v$_520_out0 };
assign v$_338_out0 = v$_658_out1[0:0];
assign v$_338_out1 = v$_658_out1[9:9];
assign v$G6_593_out0 = v$_645_out0 && v$_658_out0;
assign v$_344_out0 = { v$G5_83_out0,v$G6_593_out0 };
assign v$G7_503_out0 = v$_690_out0 && v$_338_out0;
assign v$_591_out0 = v$_338_out1[0:0];
assign v$_591_out1 = v$_338_out1[8:8];
assign v$_354_out0 = v$_591_out1[0:0];
assign v$_354_out1 = v$_591_out1[7:7];
assign v$G8_368_out0 = v$_303_out0 && v$_591_out0;
assign v$G9_167_out0 = v$_574_out0 && v$_354_out0;
assign v$_205_out0 = { v$G7_503_out0,v$G8_368_out0 };
assign v$_633_out0 = v$_354_out1[0:0];
assign v$_633_out1 = v$_354_out1[6:6];
assign v$_24_out0 = v$_633_out1[0:0];
assign v$_24_out1 = v$_633_out1[5:5];
assign v$_48_out0 = { v$_344_out0,v$_205_out0 };
assign v$G10_371_out0 = v$_346_out0 && v$_633_out0;
assign v$_85_out0 = { v$_331_out0,v$_48_out0 };
assign v$G11_159_out0 = v$_683_out0 && v$_24_out0;
assign v$_332_out0 = v$_24_out1[0:0];
assign v$_332_out1 = v$_24_out1[4:4];
assign v$_579_out0 = { v$G9_167_out0,v$G10_371_out0 };
assign v$_378_out0 = v$_332_out1[0:0];
assign v$_378_out1 = v$_332_out1[3:3];
assign v$G12_424_out0 = v$_155_out0 && v$_332_out0;
assign v$_88_out0 = v$_378_out1[0:0];
assign v$_88_out1 = v$_378_out1[2:2];
assign v$G13_246_out0 = v$_654_out0 && v$_378_out0;
assign v$_680_out0 = { v$G11_159_out0,v$G12_424_out0 };
assign v$G14_32_out0 = v$_21_out0 && v$_88_out0;
assign v$_478_out0 = { v$_579_out0,v$_680_out0 };
assign v$_709_out0 = v$_88_out1[0:0];
assign v$_709_out1 = v$_88_out1[1:1];
assign v$G16_223_out0 = v$_175_out1 && v$_709_out1;
assign v$G15_291_out0 = v$_175_out0 && v$_709_out0;
assign v$_473_out0 = { v$G13_246_out0,v$G14_32_out0 };
assign v$_463_out0 = { v$G15_291_out0,v$G16_223_out0 };
assign v$_727_out0 = { v$_473_out0,v$_463_out0 };
assign v$_528_out0 = { v$_478_out0,v$_727_out0 };
assign v$_408_out0 = { v$_85_out0,v$_528_out0 };
assign v$X_617_out0 = v$_408_out0;
assign v$ANDOUT_460_out0 = v$X_617_out0;
assign v$MUX6_91_out0 = v$G12_719_out0 ? v$ANDOUT_460_out0 : v$MUX4_725_out0;
assign v$ALUOUT_214_out0 = v$MUX6_91_out0;
assign v$ALUOUT_61_out0 = v$ALUOUT_214_out0;
assign v$MUX1_475_out0 = v$IR15_36_out0 ? v$ALUOUT_61_out0 : v$REGDIN_238_out0;
assign v$ALUOUT_477_out0 = v$ALUOUT_61_out0;
assign v$ALUOUT_506_out0 = v$ALUOUT_61_out0;
assign v$ALUOUT_174_out0 = v$ALUOUT_477_out0;
assign v$DIN3_518_out0 = v$MUX1_475_out0;
assign v$ALUOUT_721_out0 = v$ALUOUT_506_out0;
assign v$MUX12_15_out0 = v$RET_252_out0 ? v$R1S_29_out0 : v$DIN3_518_out0;
assign v$MUX11_165_out0 = v$RET_252_out0 ? v$R0S_140_out0 : v$DIN3_518_out0;
assign v$MUX14_198_out0 = v$RET_252_out0 ? v$R3S_650_out0 : v$DIN3_518_out0;
assign v$MUX13_548_out0 = v$RET_252_out0 ? v$R2S_161_out0 : v$DIN3_518_out0;


endmodule
